ram(0) <= "0110000000000000";
ram(1) <= "0010000001101001";
ram(2) <= "0110000000000000";
ram(3) <= "0010000001101000";
ram(4) <= "1000000000001000";
ram(5) <= "0001000001100100";
ram(6) <= "0110000000000001";
ram(7) <= "1001000000000000";
ram(8) <= "0001000001101000";
ram(9) <= "0100000001101001";
ram(10) <= "1000000000010001";
ram(11) <= "0001000001101001";
ram(12) <= "0010000001100111";
ram(13) <= "0001000001101000";
ram(14) <= "0010000001101001";
ram(15) <= "0001000001100111";
ram(16) <= "0010000001101000";
ram(17) <= "0001000001101001";
ram(18) <= "0010000001100110";
ram(19) <= "0001000001101001";
ram(20) <= "0010000001100100";
ram(21) <= "0001000001100110";
ram(22) <= "0100000001101010";
ram(23) <= "0111000000011010";
ram(24) <= "1000000000011010";
ram(25) <= "1001000000000101";
ram(26) <= "0001000001101001";
ram(27) <= "1110000001101000";
ram(28) <= "0010000001100101";
ram(29) <= "0001000001100101";
ram(30) <= "0111000000000101";
ram(31) <= "0010000001100100";
ram(32) <= "0001000001101000";
ram(33) <= "0010000001101001";
ram(34) <= "0001000001100101";
ram(35) <= "0010000001101000";
ram(36) <= "0001000001101010";
ram(37) <= "1100000000000001";
ram(38) <= "0010000001101010";
ram(39) <= "1001000000010101";
ram(40) <= "0000000000000000";
ram(41) <= "0000000000000000";
ram(42) <= "0000000000000000";
ram(43) <= "0000000000000000";
ram(44) <= "0000000000000000";
ram(45) <= "0000000000000000";
ram(46) <= "0000000000000000";
ram(47) <= "0000000000000000";
ram(48) <= "0000000000000000";
ram(49) <= "0000000000000000";
ram(50) <= "0000000000000000";
ram(51) <= "0000000000000000";
ram(52) <= "0000000000000000";
ram(53) <= "0000000000000000";
ram(54) <= "0000000000000000";
ram(55) <= "0000000000000000";
ram(56) <= "0000000000000000";
ram(57) <= "0000000000000000";
ram(58) <= "0000000000000000";
ram(59) <= "0000000000000000";
ram(60) <= "0000000000000000";
ram(61) <= "0000000000000000";
ram(62) <= "0000000000000000";
ram(63) <= "0000000000000000";
ram(64) <= "0000000000000000";
ram(65) <= "0000000000000000";
ram(66) <= "0000000000000000";
ram(67) <= "0000000000000000";
ram(68) <= "0000000000000000";
ram(69) <= "0000000000000000";
ram(70) <= "0000000000000000";
ram(71) <= "0000000000000000";
ram(72) <= "0000000000000000";
ram(73) <= "0000000000000000";
ram(74) <= "0000000000000000";
ram(75) <= "0000000000000000";
ram(76) <= "0000000000000000";
ram(77) <= "0000000000000000";
ram(78) <= "0000000000000000";
ram(79) <= "0000000000000000";
ram(80) <= "0000000000000000";
ram(81) <= "0000000000000000";
ram(82) <= "0000000000000000";
ram(83) <= "0000000000000000";
ram(84) <= "0000000000000000";
ram(85) <= "0000000000000000";
ram(86) <= "0000000000000000";
ram(87) <= "0000000000000000";
ram(88) <= "0000000000000000";
ram(89) <= "0000000000000000";
ram(90) <= "0000000000000000";
ram(91) <= "0000000000000000";
ram(92) <= "0000000000000000";
ram(93) <= "0000000000000000";
ram(94) <= "0000000000000000";
ram(95) <= "0000000000000000";
ram(96) <= "0000000000000000";
ram(97) <= "0000000000000000";
ram(98) <= "0000000000000000";
ram(99) <= "0000000000000000";
ram(100) <= "0000000000000000";
ram(101) <= "0000000000000000";
ram(102) <= "0000000000000000";
ram(103) <= "0000000000000000";
ram(104) <= "0000000000000000";
ram(105) <= "0000000000000000";
ram(106) <= "0000000000000000";
ram(107) <= "0000000000000000";
ram(108) <= "0000000000000000";
ram(109) <= "0000000000000000";
ram(110) <= "0000000000000000";
ram(111) <= "0000000000000000";
ram(112) <= "0000000000000000";
ram(113) <= "0000000000000000";
ram(114) <= "0000000000000000";
ram(115) <= "0000000000000000";
ram(116) <= "0000000000000000";
ram(117) <= "0000000000000000";
ram(118) <= "0000000000000000";
ram(119) <= "0000000000000000";
ram(120) <= "0000000000000000";
ram(121) <= "0000000000000000";
ram(122) <= "0000000000000000";
ram(123) <= "0000000000000000";
ram(124) <= "0000000000000000";
ram(125) <= "0000000000000000";
ram(126) <= "0000000000000000";
ram(127) <= "0000000000000000";
ram(128) <= "0000000000000000";
ram(129) <= "0000000000000000";
ram(130) <= "0000000000000000";
ram(131) <= "0000000000000000";
ram(132) <= "0000000000000000";
ram(133) <= "0000000000000000";
ram(134) <= "0000000000000000";
ram(135) <= "0000000000000000";
ram(136) <= "0000000000000000";
ram(137) <= "0000000000000000";
ram(138) <= "0000000000000000";
ram(139) <= "0000000000000000";
ram(140) <= "0000000000000000";
ram(141) <= "0000000000000000";
ram(142) <= "0000000000000000";
ram(143) <= "0000000000000000";
ram(144) <= "0000000000000000";
ram(145) <= "0000000000000000";
ram(146) <= "0000000000000000";
ram(147) <= "0000000000000000";
ram(148) <= "0000000000000000";
ram(149) <= "0000000000000000";
ram(150) <= "0000000000000000";
ram(151) <= "0000000000000000";
ram(152) <= "0000000000000000";
ram(153) <= "0000000000000000";
ram(154) <= "0000000000000000";
ram(155) <= "0000000000000000";
ram(156) <= "0000000000000000";
ram(157) <= "0000000000000000";
ram(158) <= "0000000000000000";
ram(159) <= "0000000000000000";
ram(160) <= "0000000000000000";
ram(161) <= "0000000000000000";
ram(162) <= "0000000000000000";
ram(163) <= "0000000000000000";
ram(164) <= "0000000000000000";
ram(165) <= "0000000000000000";
ram(166) <= "0000000000000000";
ram(167) <= "0000000000000000";
ram(168) <= "0000000000000000";
ram(169) <= "0000000000000000";
ram(170) <= "0000000000000000";
ram(171) <= "0000000000000000";
ram(172) <= "0000000000000000";
ram(173) <= "0000000000000000";
ram(174) <= "0000000000000000";
ram(175) <= "0000000000000000";
ram(176) <= "0000000000000000";
ram(177) <= "0000000000000000";
ram(178) <= "0000000000000000";
ram(179) <= "0000000000000000";
ram(180) <= "0000000000000000";
ram(181) <= "0000000000000000";
ram(182) <= "0000000000000000";
ram(183) <= "0000000000000000";
ram(184) <= "0000000000000000";
ram(185) <= "0000000000000000";
ram(186) <= "0000000000000000";
ram(187) <= "0000000000000000";
ram(188) <= "0000000000000000";
ram(189) <= "0000000000000000";
ram(190) <= "0000000000000000";
ram(191) <= "0000000000000000";
ram(192) <= "0000000000000000";
ram(193) <= "0000000000000000";
ram(194) <= "0000000000000000";
ram(195) <= "0000000000000000";
ram(196) <= "0000000000000000";
ram(197) <= "0000000000000000";
ram(198) <= "0000000000000000";
ram(199) <= "0000000000000000";
ram(200) <= "0000000000000000";
ram(201) <= "0000000000000000";
ram(202) <= "0000000000000000";
ram(203) <= "0000000000000000";
ram(204) <= "0000000000000000";
ram(205) <= "0000000000000000";
ram(206) <= "0000000000000000";
ram(207) <= "0000000000000000";
ram(208) <= "0000000000000000";
ram(209) <= "0000000000000000";
ram(210) <= "0000000000000000";
ram(211) <= "0000000000000000";
ram(212) <= "0000000000000000";
ram(213) <= "0000000000000000";
ram(214) <= "0000000000000000";
ram(215) <= "0000000000000000";
ram(216) <= "0000000000000000";
ram(217) <= "0000000000000000";
ram(218) <= "0000000000000000";
ram(219) <= "0000000000000000";
ram(220) <= "0000000000000000";
ram(221) <= "0000000000000000";
ram(222) <= "0000000000000000";
ram(223) <= "0000000000000000";
ram(224) <= "0000000000000000";
ram(225) <= "0000000000000000";
ram(226) <= "0000000000000000";
ram(227) <= "0000000000000000";
ram(228) <= "0000000000000000";
ram(229) <= "0000000000000000";
ram(230) <= "0000000000000000";
ram(231) <= "0000000000000000";
ram(232) <= "0000000000000000";
ram(233) <= "0000000000000000";
ram(234) <= "0000000000000000";
ram(235) <= "0000000000000000";
ram(236) <= "0000000000000000";
ram(237) <= "0000000000000000";
ram(238) <= "0000000000000000";
ram(239) <= "0000000000000000";
ram(240) <= "0000000000000000";
ram(241) <= "0000000000000000";
ram(242) <= "0000000000000000";
ram(243) <= "0000000000000000";
ram(244) <= "0000000000000000";
ram(245) <= "0000000000000000";
ram(246) <= "0000000000000000";
ram(247) <= "0000000000000000";
ram(248) <= "0000000000000000";
ram(249) <= "0000000000000000";
ram(250) <= "0000000000000000";
ram(251) <= "0000000000000000";
ram(252) <= "0000000000000000";
ram(253) <= "0000000000000000";
ram(254) <= "0000000000000000";
ram(255) <= "0000000000000000";
ram(256) <= "0000000000000000";
ram(257) <= "0000000000000000";
ram(258) <= "0000000000000000";
ram(259) <= "0000000000000000";
ram(260) <= "0000000000000000";
ram(261) <= "0000000000000000";
ram(262) <= "0000000000000000";
ram(263) <= "0000000000000000";
ram(264) <= "0000000000000000";
ram(265) <= "0000000000000000";
ram(266) <= "0000000000000000";
ram(267) <= "0000000000000000";
ram(268) <= "0000000000000000";
ram(269) <= "0000000000000000";
ram(270) <= "0000000000000000";
ram(271) <= "0000000000000000";
ram(272) <= "0000000000000000";
ram(273) <= "0000000000000000";
ram(274) <= "0000000000000000";
ram(275) <= "0000000000000000";
ram(276) <= "0000000000000000";
ram(277) <= "0000000000000000";
ram(278) <= "0000000000000000";
ram(279) <= "0000000000000000";
ram(280) <= "0000000000000000";
ram(281) <= "0000000000000000";
ram(282) <= "0000000000000000";
ram(283) <= "0000000000000000";
ram(284) <= "0000000000000000";
ram(285) <= "0000000000000000";
ram(286) <= "0000000000000000";
ram(287) <= "0000000000000000";
ram(288) <= "0000000000000000";
ram(289) <= "0000000000000000";
ram(290) <= "0000000000000000";
ram(291) <= "0000000000000000";
ram(292) <= "0000000000000000";
ram(293) <= "0000000000000000";
ram(294) <= "0000000000000000";
ram(295) <= "0000000000000000";
ram(296) <= "0000000000000000";
ram(297) <= "0000000000000000";
ram(298) <= "0000000000000000";
ram(299) <= "0000000000000000";
ram(300) <= "0000000000000000";
ram(301) <= "0000000000000000";
ram(302) <= "0000000000000000";
ram(303) <= "0000000000000000";
ram(304) <= "0000000000000000";
ram(305) <= "0000000000000000";
ram(306) <= "0000000000000000";
ram(307) <= "0000000000000000";
ram(308) <= "0000000000000000";
ram(309) <= "0000000000000000";
ram(310) <= "0000000000000000";
ram(311) <= "0000000000000000";
ram(312) <= "0000000000000000";
ram(313) <= "0000000000000000";
ram(314) <= "0000000000000000";
ram(315) <= "0000000000000000";
ram(316) <= "0000000000000000";
ram(317) <= "0000000000000000";
ram(318) <= "0000000000000000";
ram(319) <= "0000000000000000";
ram(320) <= "0000000000000000";
ram(321) <= "0000000000000000";
ram(322) <= "0000000000000000";
ram(323) <= "0000000000000000";
ram(324) <= "0000000000000000";
ram(325) <= "0000000000000000";
ram(326) <= "0000000000000000";
ram(327) <= "0000000000000000";
ram(328) <= "0000000000000000";
ram(329) <= "0000000000000000";
ram(330) <= "0000000000000000";
ram(331) <= "0000000000000000";
ram(332) <= "0000000000000000";
ram(333) <= "0000000000000000";
ram(334) <= "0000000000000000";
ram(335) <= "0000000000000000";
ram(336) <= "0000000000000000";
ram(337) <= "0000000000000000";
ram(338) <= "0000000000000000";
ram(339) <= "0000000000000000";
ram(340) <= "0000000000000000";
ram(341) <= "0000000000000000";
ram(342) <= "0000000000000000";
ram(343) <= "0000000000000000";
ram(344) <= "0000000000000000";
ram(345) <= "0000000000000000";
ram(346) <= "0000000000000000";
ram(347) <= "0000000000000000";
ram(348) <= "0000000000000000";
ram(349) <= "0000000000000000";
ram(350) <= "0000000000000000";
ram(351) <= "0000000000000000";
ram(352) <= "0000000000000000";
ram(353) <= "0000000000000000";
ram(354) <= "0000000000000000";
ram(355) <= "0000000000000000";
ram(356) <= "0000000000000000";
ram(357) <= "0000000000000000";
ram(358) <= "0000000000000000";
ram(359) <= "0000000000000000";
ram(360) <= "0000000000000000";
ram(361) <= "0000000000000000";
ram(362) <= "0000000000000000";
ram(363) <= "0000000000000000";
ram(364) <= "0000000000000000";
ram(365) <= "0000000000000000";
ram(366) <= "0000000000000000";
ram(367) <= "0000000000000000";
ram(368) <= "0000000000000000";
ram(369) <= "0000000000000000";
ram(370) <= "0000000000000000";
ram(371) <= "0000000000000000";
ram(372) <= "0000000000000000";
ram(373) <= "0000000000000000";
ram(374) <= "0000000000000000";
ram(375) <= "0000000000000000";
ram(376) <= "0000000000000000";
ram(377) <= "0000000000000000";
ram(378) <= "0000000000000000";
ram(379) <= "0000000000000000";
ram(380) <= "0000000000000000";
ram(381) <= "0000000000000000";
ram(382) <= "0000000000000000";
ram(383) <= "0000000000000000";
ram(384) <= "0000000000000000";
ram(385) <= "0000000000000000";
ram(386) <= "0000000000000000";
ram(387) <= "0000000000000000";
ram(388) <= "0000000000000000";
ram(389) <= "0000000000000000";
ram(390) <= "0000000000000000";
ram(391) <= "0000000000000000";
ram(392) <= "0000000000000000";
ram(393) <= "0000000000000000";
ram(394) <= "0000000000000000";
ram(395) <= "0000000000000000";
ram(396) <= "0000000000000000";
ram(397) <= "0000000000000000";
ram(398) <= "0000000000000000";
ram(399) <= "0000000000000000";
ram(400) <= "0000000000000000";
ram(401) <= "0000000000000000";
ram(402) <= "0000000000000000";
ram(403) <= "0000000000000000";
ram(404) <= "0000000000000000";
ram(405) <= "0000000000000000";
ram(406) <= "0000000000000000";
ram(407) <= "0000000000000000";
ram(408) <= "0000000000000000";
ram(409) <= "0000000000000000";
ram(410) <= "0000000000000000";
ram(411) <= "0000000000000000";
ram(412) <= "0000000000000000";
ram(413) <= "0000000000000000";
ram(414) <= "0000000000000000";
ram(415) <= "0000000000000000";
ram(416) <= "0000000000000000";
ram(417) <= "0000000000000000";
ram(418) <= "0000000000000000";
ram(419) <= "0000000000000000";
ram(420) <= "0000000000000000";
ram(421) <= "0000000000000000";
ram(422) <= "0000000000000000";
ram(423) <= "0000000000000000";
ram(424) <= "0000000000000000";
ram(425) <= "0000000000000000";
ram(426) <= "0000000000000000";
ram(427) <= "0000000000000000";
ram(428) <= "0000000000000000";
ram(429) <= "0000000000000000";
ram(430) <= "0000000000000000";
ram(431) <= "0000000000000000";
ram(432) <= "0000000000000000";
ram(433) <= "0000000000000000";
ram(434) <= "0000000000000000";
ram(435) <= "0000000000000000";
ram(436) <= "0000000000000000";
ram(437) <= "0000000000000000";
ram(438) <= "0000000000000000";
ram(439) <= "0000000000000000";
ram(440) <= "0000000000000000";
ram(441) <= "0000000000000000";
ram(442) <= "0000000000000000";
ram(443) <= "0000000000000000";
ram(444) <= "0000000000000000";
ram(445) <= "0000000000000000";
ram(446) <= "0000000000000000";
ram(447) <= "0000000000000000";
ram(448) <= "0000000000000000";
ram(449) <= "0000000000000000";
ram(450) <= "0000000000000000";
ram(451) <= "0000000000000000";
ram(452) <= "0000000000000000";
ram(453) <= "0000000000000000";
ram(454) <= "0000000000000000";
ram(455) <= "0000000000000000";
ram(456) <= "0000000000000000";
ram(457) <= "0000000000000000";
ram(458) <= "0000000000000000";
ram(459) <= "0000000000000000";
ram(460) <= "0000000000000000";
ram(461) <= "0000000000000000";
ram(462) <= "0000000000000000";
ram(463) <= "0000000000000000";
ram(464) <= "0000000000000000";
ram(465) <= "0000000000000000";
ram(466) <= "0000000000000000";
ram(467) <= "0000000000000000";
ram(468) <= "0000000000000000";
ram(469) <= "0000000000000000";
ram(470) <= "0000000000000000";
ram(471) <= "0000000000000000";
ram(472) <= "0000000000000000";
ram(473) <= "0000000000000000";
ram(474) <= "0000000000000000";
ram(475) <= "0000000000000000";
ram(476) <= "0000000000000000";
ram(477) <= "0000000000000000";
ram(478) <= "0000000000000000";
ram(479) <= "0000000000000000";
ram(480) <= "0000000000000000";
ram(481) <= "0000000000000000";
ram(482) <= "0000000000000000";
ram(483) <= "0000000000000000";
ram(484) <= "0000000000000000";
ram(485) <= "0000000000000000";
ram(486) <= "0000000000000000";
ram(487) <= "0000000000000000";
ram(488) <= "0000000000000000";
ram(489) <= "0000000000000000";
ram(490) <= "0000000000000000";
ram(491) <= "0000000000000000";
ram(492) <= "0000000000000000";
ram(493) <= "0000000000000000";
ram(494) <= "0000000000000000";
ram(495) <= "0000000000000000";
ram(496) <= "0000000000000000";
ram(497) <= "0000000000000000";
ram(498) <= "0000000000000000";
ram(499) <= "0000000000000000";
ram(500) <= "0000000000000000";
ram(501) <= "0000000000000000";
ram(502) <= "0000000000000000";
ram(503) <= "0000000000000000";
ram(504) <= "0000000000000000";
ram(505) <= "0000000000000000";
ram(506) <= "0000000000000000";
ram(507) <= "0000000000000000";
ram(508) <= "0000000000000000";
ram(509) <= "0000000000000000";
ram(510) <= "0000000000000000";
ram(511) <= "0000000000000000";
ram(512) <= "0000000000000000";
ram(513) <= "0000000000000000";
ram(514) <= "0000000000000000";
ram(515) <= "0000000000000000";
ram(516) <= "0000000000000000";
ram(517) <= "0000000000000000";
ram(518) <= "0000000000000000";
ram(519) <= "0000000000000000";
ram(520) <= "0000000000000000";
ram(521) <= "0000000000000000";
ram(522) <= "0000000000000000";
ram(523) <= "0000000000000000";
ram(524) <= "0000000000000000";
ram(525) <= "0000000000000000";
ram(526) <= "0000000000000000";
ram(527) <= "0000000000000000";
ram(528) <= "0000000000000000";
ram(529) <= "0000000000000000";
ram(530) <= "0000000000000000";
ram(531) <= "0000000000000000";
ram(532) <= "0000000000000000";
ram(533) <= "0000000000000000";
ram(534) <= "0000000000000000";
ram(535) <= "0000000000000000";
ram(536) <= "0000000000000000";
ram(537) <= "0000000000000000";
ram(538) <= "0000000000000000";
ram(539) <= "0000000000000000";
ram(540) <= "0000000000000000";
ram(541) <= "0000000000000000";
ram(542) <= "0000000000000000";
ram(543) <= "0000000000000000";
ram(544) <= "0000000000000000";
ram(545) <= "0000000000000000";
ram(546) <= "0000000000000000";
ram(547) <= "0000000000000000";
ram(548) <= "0000000000000000";
ram(549) <= "0000000000000000";
ram(550) <= "0000000000000000";
ram(551) <= "0000000000000000";
ram(552) <= "0000000000000000";
ram(553) <= "0000000000000000";
ram(554) <= "0000000000000000";
ram(555) <= "0000000000000000";
ram(556) <= "0000000000000000";
ram(557) <= "0000000000000000";
ram(558) <= "0000000000000000";
ram(559) <= "0000000000000000";
ram(560) <= "0000000000000000";
ram(561) <= "0000000000000000";
ram(562) <= "0000000000000000";
ram(563) <= "0000000000000000";
ram(564) <= "0000000000000000";
ram(565) <= "0000000000000000";
ram(566) <= "0000000000000000";
ram(567) <= "0000000000000000";
ram(568) <= "0000000000000000";
ram(569) <= "0000000000000000";
ram(570) <= "0000000000000000";
ram(571) <= "0000000000000000";
ram(572) <= "0000000000000000";
ram(573) <= "0000000000000000";
ram(574) <= "0000000000000000";
ram(575) <= "0000000000000000";
ram(576) <= "0000000000000000";
ram(577) <= "0000000000000000";
ram(578) <= "0000000000000000";
ram(579) <= "0000000000000000";
ram(580) <= "0000000000000000";
ram(581) <= "0000000000000000";
ram(582) <= "0000000000000000";
ram(583) <= "0000000000000000";
ram(584) <= "0000000000000000";
ram(585) <= "0000000000000000";
ram(586) <= "0000000000000000";
ram(587) <= "0000000000000000";
ram(588) <= "0000000000000000";
ram(589) <= "0000000000000000";
ram(590) <= "0000000000000000";
ram(591) <= "0000000000000000";
ram(592) <= "0000000000000000";
ram(593) <= "0000000000000000";
ram(594) <= "0000000000000000";
ram(595) <= "0000000000000000";
ram(596) <= "0000000000000000";
ram(597) <= "0000000000000000";
ram(598) <= "0000000000000000";
ram(599) <= "0000000000000000";
ram(600) <= "0000000000000000";
ram(601) <= "0000000000000000";
ram(602) <= "0000000000000000";
ram(603) <= "0000000000000000";
ram(604) <= "0000000000000000";
ram(605) <= "0000000000000000";
ram(606) <= "0000000000000000";
ram(607) <= "0000000000000000";
ram(608) <= "0000000000000000";
ram(609) <= "0000000000000000";
ram(610) <= "0000000000000000";
ram(611) <= "0000000000000000";
ram(612) <= "0000000000000000";
ram(613) <= "0000000000000000";
ram(614) <= "0000000000000000";
ram(615) <= "0000000000000000";
ram(616) <= "0000000000000000";
ram(617) <= "0000000000000000";
ram(618) <= "0000000000000000";
ram(619) <= "0000000000000000";
ram(620) <= "0000000000000000";
ram(621) <= "0000000000000000";
ram(622) <= "0000000000000000";
ram(623) <= "0000000000000000";
ram(624) <= "0000000000000000";
ram(625) <= "0000000000000000";
ram(626) <= "0000000000000000";
ram(627) <= "0000000000000000";
ram(628) <= "0000000000000000";
ram(629) <= "0000000000000000";
ram(630) <= "0000000000000000";
ram(631) <= "0000000000000000";
ram(632) <= "0000000000000000";
ram(633) <= "0000000000000000";
ram(634) <= "0000000000000000";
ram(635) <= "0000000000000000";
ram(636) <= "0000000000000000";
ram(637) <= "0000000000000000";
ram(638) <= "0000000000000000";
ram(639) <= "0000000000000000";
ram(640) <= "0000000000000000";
ram(641) <= "0000000000000000";
ram(642) <= "0000000000000000";
ram(643) <= "0000000000000000";
ram(644) <= "0000000000000000";
ram(645) <= "0000000000000000";
ram(646) <= "0000000000000000";
ram(647) <= "0000000000000000";
ram(648) <= "0000000000000000";
ram(649) <= "0000000000000000";
ram(650) <= "0000000000000000";
ram(651) <= "0000000000000000";
ram(652) <= "0000000000000000";
ram(653) <= "0000000000000000";
ram(654) <= "0000000000000000";
ram(655) <= "0000000000000000";
ram(656) <= "0000000000000000";
ram(657) <= "0000000000000000";
ram(658) <= "0000000000000000";
ram(659) <= "0000000000000000";
ram(660) <= "0000000000000000";
ram(661) <= "0000000000000000";
ram(662) <= "0000000000000000";
ram(663) <= "0000000000000000";
ram(664) <= "0000000000000000";
ram(665) <= "0000000000000000";
ram(666) <= "0000000000000000";
ram(667) <= "0000000000000000";
ram(668) <= "0000000000000000";
ram(669) <= "0000000000000000";
ram(670) <= "0000000000000000";
ram(671) <= "0000000000000000";
ram(672) <= "0000000000000000";
ram(673) <= "0000000000000000";
ram(674) <= "0000000000000000";
ram(675) <= "0000000000000000";
ram(676) <= "0000000000000000";
ram(677) <= "0000000000000000";
ram(678) <= "0000000000000000";
ram(679) <= "0000000000000000";
ram(680) <= "0000000000000000";
ram(681) <= "0000000000000000";
ram(682) <= "0000000000000000";
ram(683) <= "0000000000000000";
ram(684) <= "0000000000000000";
ram(685) <= "0000000000000000";
ram(686) <= "0000000000000000";
ram(687) <= "0000000000000000";
ram(688) <= "0000000000000000";
ram(689) <= "0000000000000000";
ram(690) <= "0000000000000000";
ram(691) <= "0000000000000000";
ram(692) <= "0000000000000000";
ram(693) <= "0000000000000000";
ram(694) <= "0000000000000000";
ram(695) <= "0000000000000000";
ram(696) <= "0000000000000000";
ram(697) <= "0000000000000000";
ram(698) <= "0000000000000000";
ram(699) <= "0000000000000000";
ram(700) <= "0000000000000000";
ram(701) <= "0000000000000000";
ram(702) <= "0000000000000000";
ram(703) <= "0000000000000000";
ram(704) <= "0000000000000000";
ram(705) <= "0000000000000000";
ram(706) <= "0000000000000000";
ram(707) <= "0000000000000000";
ram(708) <= "0000000000000000";
ram(709) <= "0000000000000000";
ram(710) <= "0000000000000000";
ram(711) <= "0000000000000000";
ram(712) <= "0000000000000000";
ram(713) <= "0000000000000000";
ram(714) <= "0000000000000000";
ram(715) <= "0000000000000000";
ram(716) <= "0000000000000000";
ram(717) <= "0000000000000000";
ram(718) <= "0000000000000000";
ram(719) <= "0000000000000000";
ram(720) <= "0000000000000000";
ram(721) <= "0000000000000000";
ram(722) <= "0000000000000000";
ram(723) <= "0000000000000000";
ram(724) <= "0000000000000000";
ram(725) <= "0000000000000000";
ram(726) <= "0000000000000000";
ram(727) <= "0000000000000000";
ram(728) <= "0000000000000000";
ram(729) <= "0000000000000000";
ram(730) <= "0000000000000000";
ram(731) <= "0000000000000000";
ram(732) <= "0000000000000000";
ram(733) <= "0000000000000000";
ram(734) <= "0000000000000000";
ram(735) <= "0000000000000000";
ram(736) <= "0000000000000000";
ram(737) <= "0000000000000000";
ram(738) <= "0000000000000000";
ram(739) <= "0000000000000000";
ram(740) <= "0000000000000000";
ram(741) <= "0000000000000000";
ram(742) <= "0000000000000000";
ram(743) <= "0000000000000000";
ram(744) <= "0000000000000000";
ram(745) <= "0000000000000000";
ram(746) <= "0000000000000000";
ram(747) <= "0000000000000000";
ram(748) <= "0000000000000000";
ram(749) <= "0000000000000000";
ram(750) <= "0000000000000000";
ram(751) <= "0000000000000000";
ram(752) <= "0000000000000000";
ram(753) <= "0000000000000000";
ram(754) <= "0000000000000000";
ram(755) <= "0000000000000000";
ram(756) <= "0000000000000000";
ram(757) <= "0000000000000000";
ram(758) <= "0000000000000000";
ram(759) <= "0000000000000000";
ram(760) <= "0000000000000000";
ram(761) <= "0000000000000000";
ram(762) <= "0000000000000000";
ram(763) <= "0000000000000000";
ram(764) <= "0000000000000000";
ram(765) <= "0000000000000000";
ram(766) <= "0000000000000000";
ram(767) <= "0000000000000000";
ram(768) <= "0000000000000000";
ram(769) <= "0000000000000000";
ram(770) <= "0000000000000000";
ram(771) <= "0000000000000000";
ram(772) <= "0000000000000000";
ram(773) <= "0000000000000000";
ram(774) <= "0000000000000000";
ram(775) <= "0000000000000000";
ram(776) <= "0000000000000000";
ram(777) <= "0000000000000000";
ram(778) <= "0000000000000000";
ram(779) <= "0000000000000000";
ram(780) <= "0000000000000000";
ram(781) <= "0000000000000000";
ram(782) <= "0000000000000000";
ram(783) <= "0000000000000000";
ram(784) <= "0000000000000000";
ram(785) <= "0000000000000000";
ram(786) <= "0000000000000000";
ram(787) <= "0000000000000000";
ram(788) <= "0000000000000000";
ram(789) <= "0000000000000000";
ram(790) <= "0000000000000000";
ram(791) <= "0000000000000000";
ram(792) <= "0000000000000000";
ram(793) <= "0000000000000000";
ram(794) <= "0000000000000000";
ram(795) <= "0000000000000000";
ram(796) <= "0000000000000000";
ram(797) <= "0000000000000000";
ram(798) <= "0000000000000000";
ram(799) <= "0000000000000000";
ram(800) <= "0000000000000000";
ram(801) <= "0000000000000000";
ram(802) <= "0000000000000000";
ram(803) <= "0000000000000000";
ram(804) <= "0000000000000000";
ram(805) <= "0000000000000000";
ram(806) <= "0000000000000000";
ram(807) <= "0000000000000000";
ram(808) <= "0000000000000000";
ram(809) <= "0000000000000000";
ram(810) <= "0000000000000000";
ram(811) <= "0000000000000000";
ram(812) <= "0000000000000000";
ram(813) <= "0000000000000000";
ram(814) <= "0000000000000000";
ram(815) <= "0000000000000000";
ram(816) <= "0000000000000000";
ram(817) <= "0000000000000000";
ram(818) <= "0000000000000000";
ram(819) <= "0000000000000000";
ram(820) <= "0000000000000000";
ram(821) <= "0000000000000000";
ram(822) <= "0000000000000000";
ram(823) <= "0000000000000000";
ram(824) <= "0000000000000000";
ram(825) <= "0000000000000000";
ram(826) <= "0000000000000000";
ram(827) <= "0000000000000000";
ram(828) <= "0000000000000000";
ram(829) <= "0000000000000000";
ram(830) <= "0000000000000000";
ram(831) <= "0000000000000000";
ram(832) <= "0000000000000000";
ram(833) <= "0000000000000000";
ram(834) <= "0000000000000000";
ram(835) <= "0000000000000000";
ram(836) <= "0000000000000000";
ram(837) <= "0000000000000000";
ram(838) <= "0000000000000000";
ram(839) <= "0000000000000000";
ram(840) <= "0000000000000000";
ram(841) <= "0000000000000000";
ram(842) <= "0000000000000000";
ram(843) <= "0000000000000000";
ram(844) <= "0000000000000000";
ram(845) <= "0000000000000000";
ram(846) <= "0000000000000000";
ram(847) <= "0000000000000000";
ram(848) <= "0000000000000000";
ram(849) <= "0000000000000000";
ram(850) <= "0000000000000000";
ram(851) <= "0000000000000000";
ram(852) <= "0000000000000000";
ram(853) <= "0000000000000000";
ram(854) <= "0000000000000000";
ram(855) <= "0000000000000000";
ram(856) <= "0000000000000000";
ram(857) <= "0000000000000000";
ram(858) <= "0000000000000000";
ram(859) <= "0000000000000000";
ram(860) <= "0000000000000000";
ram(861) <= "0000000000000000";
ram(862) <= "0000000000000000";
ram(863) <= "0000000000000000";
ram(864) <= "0000000000000000";
ram(865) <= "0000000000000000";
ram(866) <= "0000000000000000";
ram(867) <= "0000000000000000";
ram(868) <= "0000000000000000";
ram(869) <= "0000000000000000";
ram(870) <= "0000000000000000";
ram(871) <= "0000000000000000";
ram(872) <= "0000000000000000";
ram(873) <= "0000000000000000";
ram(874) <= "0000000000000000";
ram(875) <= "0000000000000000";
ram(876) <= "0000000000000000";
ram(877) <= "0000000000000000";
ram(878) <= "0000000000000000";
ram(879) <= "0000000000000000";
ram(880) <= "0000000000000000";
ram(881) <= "0000000000000000";
ram(882) <= "0000000000000000";
ram(883) <= "0000000000000000";
ram(884) <= "0000000000000000";
ram(885) <= "0000000000000000";
ram(886) <= "0000000000000000";
ram(887) <= "0000000000000000";
ram(888) <= "0000000000000000";
ram(889) <= "0000000000000000";
ram(890) <= "0000000000000000";
ram(891) <= "0000000000000000";
ram(892) <= "0000000000000000";
ram(893) <= "0000000000000000";
ram(894) <= "0000000000000000";
ram(895) <= "0000000000000000";
ram(896) <= "0000000000000000";
ram(897) <= "0000000000000000";
ram(898) <= "0000000000000000";
ram(899) <= "0000000000000000";
ram(900) <= "0000000000000000";
ram(901) <= "0000000000000000";
ram(902) <= "0000000000000000";
ram(903) <= "0000000000000000";
ram(904) <= "0000000000000000";
ram(905) <= "0000000000000000";
ram(906) <= "0000000000000000";
ram(907) <= "0000000000000000";
ram(908) <= "0000000000000000";
ram(909) <= "0000000000000000";
ram(910) <= "0000000000000000";
ram(911) <= "0000000000000000";
ram(912) <= "0000000000000000";
ram(913) <= "0000000000000000";
ram(914) <= "0000000000000000";
ram(915) <= "0000000000000000";
ram(916) <= "0000000000000000";
ram(917) <= "0000000000000000";
ram(918) <= "0000000000000000";
ram(919) <= "0000000000000000";
ram(920) <= "0000000000000000";
ram(921) <= "0000000000000000";
ram(922) <= "0000000000000000";
ram(923) <= "0000000000000000";
ram(924) <= "0000000000000000";
ram(925) <= "0000000000000000";
ram(926) <= "0000000000000000";
ram(927) <= "0000000000000000";
ram(928) <= "0000000000000000";
ram(929) <= "0000000000000000";
ram(930) <= "0000000000000000";
ram(931) <= "0000000000000000";
ram(932) <= "0000000000000000";
ram(933) <= "0000000000000000";
ram(934) <= "0000000000000000";
ram(935) <= "0000000000000000";
ram(936) <= "0000000000000000";
ram(937) <= "0000000000000000";
ram(938) <= "0000000000000000";
ram(939) <= "0000000000000000";
ram(940) <= "0000000000000000";
ram(941) <= "0000000000000000";
ram(942) <= "0000000000000000";
ram(943) <= "0000000000000000";
ram(944) <= "0000000000000000";
ram(945) <= "0000000000000000";
ram(946) <= "0000000000000000";
ram(947) <= "0000000000000000";
ram(948) <= "0000000000000000";
ram(949) <= "0000000000000000";
ram(950) <= "0000000000000000";
ram(951) <= "0000000000000000";
ram(952) <= "0000000000000000";
ram(953) <= "0000000000000000";
ram(954) <= "0000000000000000";
ram(955) <= "0000000000000000";
ram(956) <= "0000000000000000";
ram(957) <= "0000000000000000";
ram(958) <= "0000000000000000";
ram(959) <= "0000000000000000";
ram(960) <= "0000000000000000";
ram(961) <= "0000000000000000";
ram(962) <= "0000000000000000";
ram(963) <= "0000000000000000";
ram(964) <= "0000000000000000";
ram(965) <= "0000000000000000";
ram(966) <= "0000000000000000";
ram(967) <= "0000000000000000";
ram(968) <= "0000000000000000";
ram(969) <= "0000000000000000";
ram(970) <= "0000000000000000";
ram(971) <= "0000000000000000";
ram(972) <= "0000000000000000";
ram(973) <= "0000000000000000";
ram(974) <= "0000000000000000";
ram(975) <= "0000000000000000";
ram(976) <= "0000000000000000";
ram(977) <= "0000000000000000";
ram(978) <= "0000000000000000";
ram(979) <= "0000000000000000";
ram(980) <= "0000000000000000";
ram(981) <= "0000000000000000";
ram(982) <= "0000000000000000";
ram(983) <= "0000000000000000";
ram(984) <= "0000000000000000";
ram(985) <= "0000000000000000";
ram(986) <= "0000000000000000";
ram(987) <= "0000000000000000";
ram(988) <= "0000000000000000";
ram(989) <= "0000000000000000";
ram(990) <= "0000000000000000";
ram(991) <= "0000000000000000";
ram(992) <= "0000000000000000";
ram(993) <= "0000000000000000";
ram(994) <= "0000000000000000";
ram(995) <= "0000000000000000";
ram(996) <= "0000000000000000";
ram(997) <= "0000000000000000";
ram(998) <= "0000000000000000";
ram(999) <= "0000000000000000";
ram(1000) <= "0000000000000000";
ram(1001) <= "0000000000000000";
ram(1002) <= "0000000000000000";
ram(1003) <= "0000000000000000";
ram(1004) <= "0000000000000000";
ram(1005) <= "0000000000000000";
ram(1006) <= "0000000000000000";
ram(1007) <= "0000000000000000";
ram(1008) <= "0000000000000000";
ram(1009) <= "0000000000000000";
ram(1010) <= "0000000000000000";
ram(1011) <= "0000000000000000";
ram(1012) <= "0000000000000000";
ram(1013) <= "0000000000000000";
ram(1014) <= "0000000000000000";
ram(1015) <= "0000000000000000";
ram(1016) <= "0000000000000000";
ram(1017) <= "0000000000000000";
ram(1018) <= "0000000000000000";
ram(1019) <= "0000000000000000";
ram(1020) <= "0000000000000000";
ram(1021) <= "0000000000000000";
ram(1022) <= "0000000000000000";
ram(1023) <= "0000000000000000";
ram(1024) <= "0000000000000000";
ram(1025) <= "0000000000000000";
ram(1026) <= "0000000000000000";
ram(1027) <= "0000000000000000";
ram(1028) <= "0000000000000000";
ram(1029) <= "0000000000000000";
ram(1030) <= "0000000000000000";
ram(1031) <= "0000000000000000";
ram(1032) <= "0000000000000000";
ram(1033) <= "0000000000000000";
ram(1034) <= "0000000000000000";
ram(1035) <= "0000000000000000";
ram(1036) <= "0000000000000000";
ram(1037) <= "0000000000000000";
ram(1038) <= "0000000000000000";
ram(1039) <= "0000000000000000";
ram(1040) <= "0000000000000000";
ram(1041) <= "0000000000000000";
ram(1042) <= "0000000000000000";
ram(1043) <= "0000000000000000";
ram(1044) <= "0000000000000000";
ram(1045) <= "0000000000000000";
ram(1046) <= "0000000000000000";
ram(1047) <= "0000000000000000";
ram(1048) <= "0000000000000000";
ram(1049) <= "0000000000000000";
ram(1050) <= "0000000000000000";
ram(1051) <= "0000000000000000";
ram(1052) <= "0000000000000000";
ram(1053) <= "0000000000000000";
ram(1054) <= "0000000000000000";
ram(1055) <= "0000000000000000";
ram(1056) <= "0000000000000000";
ram(1057) <= "0000000000000000";
ram(1058) <= "0000000000000000";
ram(1059) <= "0000000000000000";
ram(1060) <= "0000000000000000";
ram(1061) <= "0000000000000000";
ram(1062) <= "0000000000000000";
ram(1063) <= "0000000000000000";
ram(1064) <= "0000000000000000";
ram(1065) <= "0000000000000000";
ram(1066) <= "0000000000000000";
ram(1067) <= "0000000000000000";
ram(1068) <= "0000000000000000";
ram(1069) <= "0000000000000000";
ram(1070) <= "0000000000000000";
ram(1071) <= "0000000000000000";
ram(1072) <= "0000000000000000";
ram(1073) <= "0000000000000000";
ram(1074) <= "0000000000000000";
ram(1075) <= "0000000000000000";
ram(1076) <= "0000000000000000";
ram(1077) <= "0000000000000000";
ram(1078) <= "0000000000000000";
ram(1079) <= "0000000000000000";
ram(1080) <= "0000000000000000";
ram(1081) <= "0000000000000000";
ram(1082) <= "0000000000000000";
ram(1083) <= "0000000000000000";
ram(1084) <= "0000000000000000";
ram(1085) <= "0000000000000000";
ram(1086) <= "0000000000000000";
ram(1087) <= "0000000000000000";
ram(1088) <= "0000000000000000";
ram(1089) <= "0000000000000000";
ram(1090) <= "0000000000000000";
ram(1091) <= "0000000000000000";
ram(1092) <= "0000000000000000";
ram(1093) <= "0000000000000000";
ram(1094) <= "0000000000000000";
ram(1095) <= "0000000000000000";
ram(1096) <= "0000000000000000";
ram(1097) <= "0000000000000000";
ram(1098) <= "0000000000000000";
ram(1099) <= "0000000000000000";
ram(1100) <= "0000000000000000";
ram(1101) <= "0000000000000000";
ram(1102) <= "0000000000000000";
ram(1103) <= "0000000000000000";
ram(1104) <= "0000000000000000";
ram(1105) <= "0000000000000000";
ram(1106) <= "0000000000000000";
ram(1107) <= "0000000000000000";
ram(1108) <= "0000000000000000";
ram(1109) <= "0000000000000000";
ram(1110) <= "0000000000000000";
ram(1111) <= "0000000000000000";
ram(1112) <= "0000000000000000";
ram(1113) <= "0000000000000000";
ram(1114) <= "0000000000000000";
ram(1115) <= "0000000000000000";
ram(1116) <= "0000000000000000";
ram(1117) <= "0000000000000000";
ram(1118) <= "0000000000000000";
ram(1119) <= "0000000000000000";
ram(1120) <= "0000000000000000";
ram(1121) <= "0000000000000000";
ram(1122) <= "0000000000000000";
ram(1123) <= "0000000000000000";
ram(1124) <= "0000000000000000";
ram(1125) <= "0000000000000000";
ram(1126) <= "0000000000000000";
ram(1127) <= "0000000000000000";
ram(1128) <= "0000000000000000";
ram(1129) <= "0000000000000000";
ram(1130) <= "0000000000000000";
ram(1131) <= "0000000000000000";
ram(1132) <= "0000000000000000";
ram(1133) <= "0000000000000000";
ram(1134) <= "0000000000000000";
ram(1135) <= "0000000000000000";
ram(1136) <= "0000000000000000";
ram(1137) <= "0000000000000000";
ram(1138) <= "0000000000000000";
ram(1139) <= "0000000000000000";
ram(1140) <= "0000000000000000";
ram(1141) <= "0000000000000000";
ram(1142) <= "0000000000000000";
ram(1143) <= "0000000000000000";
ram(1144) <= "0000000000000000";
ram(1145) <= "0000000000000000";
ram(1146) <= "0000000000000000";
ram(1147) <= "0000000000000000";
ram(1148) <= "0000000000000000";
ram(1149) <= "0000000000000000";
ram(1150) <= "0000000000000000";
ram(1151) <= "0000000000000000";
ram(1152) <= "0000000000000000";
ram(1153) <= "0000000000000000";
ram(1154) <= "0000000000000000";
ram(1155) <= "0000000000000000";
ram(1156) <= "0000000000000000";
ram(1157) <= "0000000000000000";
ram(1158) <= "0000000000000000";
ram(1159) <= "0000000000000000";
ram(1160) <= "0000000000000000";
ram(1161) <= "0000000000000000";
ram(1162) <= "0000000000000000";
ram(1163) <= "0000000000000000";
ram(1164) <= "0000000000000000";
ram(1165) <= "0000000000000000";
ram(1166) <= "0000000000000000";
ram(1167) <= "0000000000000000";
ram(1168) <= "0000000000000000";
ram(1169) <= "0000000000000000";
ram(1170) <= "0000000000000000";
ram(1171) <= "0000000000000000";
ram(1172) <= "0000000000000000";
ram(1173) <= "0000000000000000";
ram(1174) <= "0000000000000000";
ram(1175) <= "0000000000000000";
ram(1176) <= "0000000000000000";
ram(1177) <= "0000000000000000";
ram(1178) <= "0000000000000000";
ram(1179) <= "0000000000000000";
ram(1180) <= "0000000000000000";
ram(1181) <= "0000000000000000";
ram(1182) <= "0000000000000000";
ram(1183) <= "0000000000000000";
ram(1184) <= "0000000000000000";
ram(1185) <= "0000000000000000";
ram(1186) <= "0000000000000000";
ram(1187) <= "0000000000000000";
ram(1188) <= "0000000000000000";
ram(1189) <= "0000000000000000";
ram(1190) <= "0000000000000000";
ram(1191) <= "0000000000000000";
ram(1192) <= "0000000000000000";
ram(1193) <= "0000000000000000";
ram(1194) <= "0000000000000000";
ram(1195) <= "0000000000000000";
ram(1196) <= "0000000000000000";
ram(1197) <= "0000000000000000";
ram(1198) <= "0000000000000000";
ram(1199) <= "0000000000000000";
ram(1200) <= "0000000000000000";
ram(1201) <= "0000000000000000";
ram(1202) <= "0000000000000000";
ram(1203) <= "0000000000000000";
ram(1204) <= "0000000000000000";
ram(1205) <= "0000000000000000";
ram(1206) <= "0000000000000000";
ram(1207) <= "0000000000000000";
ram(1208) <= "0000000000000000";
ram(1209) <= "0000000000000000";
ram(1210) <= "0000000000000000";
ram(1211) <= "0000000000000000";
ram(1212) <= "0000000000000000";
ram(1213) <= "0000000000000000";
ram(1214) <= "0000000000000000";
ram(1215) <= "0000000000000000";
ram(1216) <= "0000000000000000";
ram(1217) <= "0000000000000000";
ram(1218) <= "0000000000000000";
ram(1219) <= "0000000000000000";
ram(1220) <= "0000000000000000";
ram(1221) <= "0000000000000000";
ram(1222) <= "0000000000000000";
ram(1223) <= "0000000000000000";
ram(1224) <= "0000000000000000";
ram(1225) <= "0000000000000000";
ram(1226) <= "0000000000000000";
ram(1227) <= "0000000000000000";
ram(1228) <= "0000000000000000";
ram(1229) <= "0000000000000000";
ram(1230) <= "0000000000000000";
ram(1231) <= "0000000000000000";
ram(1232) <= "0000000000000000";
ram(1233) <= "0000000000000000";
ram(1234) <= "0000000000000000";
ram(1235) <= "0000000000000000";
ram(1236) <= "0000000000000000";
ram(1237) <= "0000000000000000";
ram(1238) <= "0000000000000000";
ram(1239) <= "0000000000000000";
ram(1240) <= "0000000000000000";
ram(1241) <= "0000000000000000";
ram(1242) <= "0000000000000000";
ram(1243) <= "0000000000000000";
ram(1244) <= "0000000000000000";
ram(1245) <= "0000000000000000";
ram(1246) <= "0000000000000000";
ram(1247) <= "0000000000000000";
ram(1248) <= "0000000000000000";
ram(1249) <= "0000000000000000";
ram(1250) <= "0000000000000000";
ram(1251) <= "0000000000000000";
ram(1252) <= "0000000000000000";
ram(1253) <= "0000000000000000";
ram(1254) <= "0000000000000000";
ram(1255) <= "0000000000000000";
ram(1256) <= "0000000000000000";
ram(1257) <= "0000000000000000";
ram(1258) <= "0000000000000000";
ram(1259) <= "0000000000000000";
ram(1260) <= "0000000000000000";
ram(1261) <= "0000000000000000";
ram(1262) <= "0000000000000000";
ram(1263) <= "0000000000000000";
ram(1264) <= "0000000000000000";
ram(1265) <= "0000000000000000";
ram(1266) <= "0000000000000000";
ram(1267) <= "0000000000000000";
ram(1268) <= "0000000000000000";
ram(1269) <= "0000000000000000";
ram(1270) <= "0000000000000000";
ram(1271) <= "0000000000000000";
ram(1272) <= "0000000000000000";
ram(1273) <= "0000000000000000";
ram(1274) <= "0000000000000000";
ram(1275) <= "0000000000000000";
ram(1276) <= "0000000000000000";
ram(1277) <= "0000000000000000";
ram(1278) <= "0000000000000000";
ram(1279) <= "0000000000000000";
ram(1280) <= "0000000000000000";
ram(1281) <= "0000000000000000";
ram(1282) <= "0000000000000000";
ram(1283) <= "0000000000000000";
ram(1284) <= "0000000000000000";
ram(1285) <= "0000000000000000";
ram(1286) <= "0000000000000000";
ram(1287) <= "0000000000000000";
ram(1288) <= "0000000000000000";
ram(1289) <= "0000000000000000";
ram(1290) <= "0000000000000000";
ram(1291) <= "0000000000000000";
ram(1292) <= "0000000000000000";
ram(1293) <= "0000000000000000";
ram(1294) <= "0000000000000000";
ram(1295) <= "0000000000000000";
ram(1296) <= "0000000000000000";
ram(1297) <= "0000000000000000";
ram(1298) <= "0000000000000000";
ram(1299) <= "0000000000000000";
ram(1300) <= "0000000000000000";
ram(1301) <= "0000000000000000";
ram(1302) <= "0000000000000000";
ram(1303) <= "0000000000000000";
ram(1304) <= "0000000000000000";
ram(1305) <= "0000000000000000";
ram(1306) <= "0000000000000000";
ram(1307) <= "0000000000000000";
ram(1308) <= "0000000000000000";
ram(1309) <= "0000000000000000";
ram(1310) <= "0000000000000000";
ram(1311) <= "0000000000000000";
ram(1312) <= "0000000000000000";
ram(1313) <= "0000000000000000";
ram(1314) <= "0000000000000000";
ram(1315) <= "0000000000000000";
ram(1316) <= "0000000000000000";
ram(1317) <= "0000000000000000";
ram(1318) <= "0000000000000000";
ram(1319) <= "0000000000000000";
ram(1320) <= "0000000000000000";
ram(1321) <= "0000000000000000";
ram(1322) <= "0000000000000000";
ram(1323) <= "0000000000000000";
ram(1324) <= "0000000000000000";
ram(1325) <= "0000000000000000";
ram(1326) <= "0000000000000000";
ram(1327) <= "0000000000000000";
ram(1328) <= "0000000000000000";
ram(1329) <= "0000000000000000";
ram(1330) <= "0000000000000000";
ram(1331) <= "0000000000000000";
ram(1332) <= "0000000000000000";
ram(1333) <= "0000000000000000";
ram(1334) <= "0000000000000000";
ram(1335) <= "0000000000000000";
ram(1336) <= "0000000000000000";
ram(1337) <= "0000000000000000";
ram(1338) <= "0000000000000000";
ram(1339) <= "0000000000000000";
ram(1340) <= "0000000000000000";
ram(1341) <= "0000000000000000";
ram(1342) <= "0000000000000000";
ram(1343) <= "0000000000000000";
ram(1344) <= "0000000000000000";
ram(1345) <= "0000000000000000";
ram(1346) <= "0000000000000000";
ram(1347) <= "0000000000000000";
ram(1348) <= "0000000000000000";
ram(1349) <= "0000000000000000";
ram(1350) <= "0000000000000000";
ram(1351) <= "0000000000000000";
ram(1352) <= "0000000000000000";
ram(1353) <= "0000000000000000";
ram(1354) <= "0000000000000000";
ram(1355) <= "0000000000000000";
ram(1356) <= "0000000000000000";
ram(1357) <= "0000000000000000";
ram(1358) <= "0000000000000000";
ram(1359) <= "0000000000000000";
ram(1360) <= "0000000000000000";
ram(1361) <= "0000000000000000";
ram(1362) <= "0000000000000000";
ram(1363) <= "0000000000000000";
ram(1364) <= "0000000000000000";
ram(1365) <= "0000000000000000";
ram(1366) <= "0000000000000000";
ram(1367) <= "0000000000000000";
ram(1368) <= "0000000000000000";
ram(1369) <= "0000000000000000";
ram(1370) <= "0000000000000000";
ram(1371) <= "0000000000000000";
ram(1372) <= "0000000000000000";
ram(1373) <= "0000000000000000";
ram(1374) <= "0000000000000000";
ram(1375) <= "0000000000000000";
ram(1376) <= "0000000000000000";
ram(1377) <= "0000000000000000";
ram(1378) <= "0000000000000000";
ram(1379) <= "0000000000000000";
ram(1380) <= "0000000000000000";
ram(1381) <= "0000000000000000";
ram(1382) <= "0000000000000000";
ram(1383) <= "0000000000000000";
ram(1384) <= "0000000000000000";
ram(1385) <= "0000000000000000";
ram(1386) <= "0000000000000000";
ram(1387) <= "0000000000000000";
ram(1388) <= "0000000000000000";
ram(1389) <= "0000000000000000";
ram(1390) <= "0000000000000000";
ram(1391) <= "0000000000000000";
ram(1392) <= "0000000000000000";
ram(1393) <= "0000000000000000";
ram(1394) <= "0000000000000000";
ram(1395) <= "0000000000000000";
ram(1396) <= "0000000000000000";
ram(1397) <= "0000000000000000";
ram(1398) <= "0000000000000000";
ram(1399) <= "0000000000000000";
ram(1400) <= "0000000000000000";
ram(1401) <= "0000000000000000";
ram(1402) <= "0000000000000000";
ram(1403) <= "0000000000000000";
ram(1404) <= "0000000000000000";
ram(1405) <= "0000000000000000";
ram(1406) <= "0000000000000000";
ram(1407) <= "0000000000000000";
ram(1408) <= "0000000000000000";
ram(1409) <= "0000000000000000";
ram(1410) <= "0000000000000000";
ram(1411) <= "0000000000000000";
ram(1412) <= "0000000000000000";
ram(1413) <= "0000000000000000";
ram(1414) <= "0000000000000000";
ram(1415) <= "0000000000000000";
ram(1416) <= "0000000000000000";
ram(1417) <= "0000000000000000";
ram(1418) <= "0000000000000000";
ram(1419) <= "0000000000000000";
ram(1420) <= "0000000000000000";
ram(1421) <= "0000000000000000";
ram(1422) <= "0000000000000000";
ram(1423) <= "0000000000000000";
ram(1424) <= "0000000000000000";
ram(1425) <= "0000000000000000";
ram(1426) <= "0000000000000000";
ram(1427) <= "0000000000000000";
ram(1428) <= "0000000000000000";
ram(1429) <= "0000000000000000";
ram(1430) <= "0000000000000000";
ram(1431) <= "0000000000000000";
ram(1432) <= "0000000000000000";
ram(1433) <= "0000000000000000";
ram(1434) <= "0000000000000000";
ram(1435) <= "0000000000000000";
ram(1436) <= "0000000000000000";
ram(1437) <= "0000000000000000";
ram(1438) <= "0000000000000000";
ram(1439) <= "0000000000000000";
ram(1440) <= "0000000000000000";
ram(1441) <= "0000000000000000";
ram(1442) <= "0000000000000000";
ram(1443) <= "0000000000000000";
ram(1444) <= "0000000000000000";
ram(1445) <= "0000000000000000";
ram(1446) <= "0000000000000000";
ram(1447) <= "0000000000000000";
ram(1448) <= "0000000000000000";
ram(1449) <= "0000000000000000";
ram(1450) <= "0000000000000000";
ram(1451) <= "0000000000000000";
ram(1452) <= "0000000000000000";
ram(1453) <= "0000000000000000";
ram(1454) <= "0000000000000000";
ram(1455) <= "0000000000000000";
ram(1456) <= "0000000000000000";
ram(1457) <= "0000000000000000";
ram(1458) <= "0000000000000000";
ram(1459) <= "0000000000000000";
ram(1460) <= "0000000000000000";
ram(1461) <= "0000000000000000";
ram(1462) <= "0000000000000000";
ram(1463) <= "0000000000000000";
ram(1464) <= "0000000000000000";
ram(1465) <= "0000000000000000";
ram(1466) <= "0000000000000000";
ram(1467) <= "0000000000000000";
ram(1468) <= "0000000000000000";
ram(1469) <= "0000000000000000";
ram(1470) <= "0000000000000000";
ram(1471) <= "0000000000000000";
ram(1472) <= "0000000000000000";
ram(1473) <= "0000000000000000";
ram(1474) <= "0000000000000000";
ram(1475) <= "0000000000000000";
ram(1476) <= "0000000000000000";
ram(1477) <= "0000000000000000";
ram(1478) <= "0000000000000000";
ram(1479) <= "0000000000000000";
ram(1480) <= "0000000000000000";
ram(1481) <= "0000000000000000";
ram(1482) <= "0000000000000000";
ram(1483) <= "0000000000000000";
ram(1484) <= "0000000000000000";
ram(1485) <= "0000000000000000";
ram(1486) <= "0000000000000000";
ram(1487) <= "0000000000000000";
ram(1488) <= "0000000000000000";
ram(1489) <= "0000000000000000";
ram(1490) <= "0000000000000000";
ram(1491) <= "0000000000000000";
ram(1492) <= "0000000000000000";
ram(1493) <= "0000000000000000";
ram(1494) <= "0000000000000000";
ram(1495) <= "0000000000000000";
ram(1496) <= "0000000000000000";
ram(1497) <= "0000000000000000";
ram(1498) <= "0000000000000000";
ram(1499) <= "0000000000000000";
ram(1500) <= "0000000000000000";
ram(1501) <= "0000000000000000";
ram(1502) <= "0000000000000000";
ram(1503) <= "0000000000000000";
ram(1504) <= "0000000000000000";
ram(1505) <= "0000000000000000";
ram(1506) <= "0000000000000000";
ram(1507) <= "0000000000000000";
ram(1508) <= "0000000000000000";
ram(1509) <= "0000000000000000";
ram(1510) <= "0000000000000000";
ram(1511) <= "0000000000000000";
ram(1512) <= "0000000000000000";
ram(1513) <= "0000000000000000";
ram(1514) <= "0000000000000000";
ram(1515) <= "0000000000000000";
ram(1516) <= "0000000000000000";
ram(1517) <= "0000000000000000";
ram(1518) <= "0000000000000000";
ram(1519) <= "0000000000000000";
ram(1520) <= "0000000000000000";
ram(1521) <= "0000000000000000";
ram(1522) <= "0000000000000000";
ram(1523) <= "0000000000000000";
ram(1524) <= "0000000000000000";
ram(1525) <= "0000000000000000";
ram(1526) <= "0000000000000000";
ram(1527) <= "0000000000000000";
ram(1528) <= "0000000000000000";
ram(1529) <= "0000000000000000";
ram(1530) <= "0000000000000000";
ram(1531) <= "0000000000000000";
ram(1532) <= "0000000000000000";
ram(1533) <= "0000000000000000";
ram(1534) <= "0000000000000000";
ram(1535) <= "0000000000000000";
ram(1536) <= "0000000000000000";
ram(1537) <= "0000000000000000";
ram(1538) <= "0000000000000000";
ram(1539) <= "0000000000000000";
ram(1540) <= "0000000000000000";
ram(1541) <= "0000000000000000";
ram(1542) <= "0000000000000000";
ram(1543) <= "0000000000000000";
ram(1544) <= "0000000000000000";
ram(1545) <= "0000000000000000";
ram(1546) <= "0000000000000000";
ram(1547) <= "0000000000000000";
ram(1548) <= "0000000000000000";
ram(1549) <= "0000000000000000";
ram(1550) <= "0000000000000000";
ram(1551) <= "0000000000000000";
ram(1552) <= "0000000000000000";
ram(1553) <= "0000000000000000";
ram(1554) <= "0000000000000000";
ram(1555) <= "0000000000000000";
ram(1556) <= "0000000000000000";
ram(1557) <= "0000000000000000";
ram(1558) <= "0000000000000000";
ram(1559) <= "0000000000000000";
ram(1560) <= "0000000000000000";
ram(1561) <= "0000000000000000";
ram(1562) <= "0000000000000000";
ram(1563) <= "0000000000000000";
ram(1564) <= "0000000000000000";
ram(1565) <= "0000000000000000";
ram(1566) <= "0000000000000000";
ram(1567) <= "0000000000000000";
ram(1568) <= "0000000000000000";
ram(1569) <= "0000000000000000";
ram(1570) <= "0000000000000000";
ram(1571) <= "0000000000000000";
ram(1572) <= "0000000000000000";
ram(1573) <= "0000000000000000";
ram(1574) <= "0000000000000000";
ram(1575) <= "0000000000000000";
ram(1576) <= "0000000000000000";
ram(1577) <= "0000000000000000";
ram(1578) <= "0000000000000000";
ram(1579) <= "0000000000000000";
ram(1580) <= "0000000000000000";
ram(1581) <= "0000000000000000";
ram(1582) <= "0000000000000000";
ram(1583) <= "0000000000000000";
ram(1584) <= "0000000000000000";
ram(1585) <= "0000000000000000";
ram(1586) <= "0000000000000000";
ram(1587) <= "0000000000000000";
ram(1588) <= "0000000000000000";
ram(1589) <= "0000000000000000";
ram(1590) <= "0000000000000000";
ram(1591) <= "0000000000000000";
ram(1592) <= "0000000000000000";
ram(1593) <= "0000000000000000";
ram(1594) <= "0000000000000000";
ram(1595) <= "0000000000000000";
ram(1596) <= "0000000000000000";
ram(1597) <= "0000000000000000";
ram(1598) <= "0000000000000000";
ram(1599) <= "0000000000000000";
ram(1600) <= "0000000000000000";
ram(1601) <= "0000000000000000";
ram(1602) <= "0000000000000000";
ram(1603) <= "0000000000000000";
ram(1604) <= "0000000000000000";
ram(1605) <= "0000000000000000";
ram(1606) <= "0000000000000000";
ram(1607) <= "0000000000000000";
ram(1608) <= "0000000000000000";
ram(1609) <= "0000000000000000";
ram(1610) <= "0000000000000000";
ram(1611) <= "0000000000000000";
ram(1612) <= "0000000000000000";
ram(1613) <= "0000000000000000";
ram(1614) <= "0000000000000000";
ram(1615) <= "0000000000000000";
ram(1616) <= "0000000000000000";
ram(1617) <= "0000000000000000";
ram(1618) <= "0000000000000000";
ram(1619) <= "0000000000000000";
ram(1620) <= "0000000000000000";
ram(1621) <= "0000000000000000";
ram(1622) <= "0000000000000000";
ram(1623) <= "0000000000000000";
ram(1624) <= "0000000000000000";
ram(1625) <= "0000000000000000";
ram(1626) <= "0000000000000000";
ram(1627) <= "0000000000000000";
ram(1628) <= "0000000000000000";
ram(1629) <= "0000000000000000";
ram(1630) <= "0000000000000000";
ram(1631) <= "0000000000000000";
ram(1632) <= "0000000000000000";
ram(1633) <= "0000000000000000";
ram(1634) <= "0000000000000000";
ram(1635) <= "0000000000000000";
ram(1636) <= "0000000000000000";
ram(1637) <= "0000000000000000";
ram(1638) <= "0000000000000000";
ram(1639) <= "0000000000000000";
ram(1640) <= "0000000000000000";
ram(1641) <= "0000000000000000";
ram(1642) <= "0000000000000000";
ram(1643) <= "0000000000000000";
ram(1644) <= "0000000000000000";
ram(1645) <= "0000000000000000";
ram(1646) <= "0000000000000000";
ram(1647) <= "0000000000000000";
ram(1648) <= "0000000000000000";
ram(1649) <= "0000000000000000";
ram(1650) <= "0000000000000000";
ram(1651) <= "0000000000000000";
ram(1652) <= "0000000000000000";
ram(1653) <= "0000000000000000";
ram(1654) <= "0000000000000000";
ram(1655) <= "0000000000000000";
ram(1656) <= "0000000000000000";
ram(1657) <= "0000000000000000";
ram(1658) <= "0000000000000000";
ram(1659) <= "0000000000000000";
ram(1660) <= "0000000000000000";
ram(1661) <= "0000000000000000";
ram(1662) <= "0000000000000000";
ram(1663) <= "0000000000000000";
ram(1664) <= "0000000000000000";
ram(1665) <= "0000000000000000";
ram(1666) <= "0000000000000000";
ram(1667) <= "0000000000000000";
ram(1668) <= "0000000000000000";
ram(1669) <= "0000000000000000";
ram(1670) <= "0000000000000000";
ram(1671) <= "0000000000000000";
ram(1672) <= "0000000000000000";
ram(1673) <= "0000000000000000";
ram(1674) <= "0000000000000000";
ram(1675) <= "0000000000000000";
ram(1676) <= "0000000000000000";
ram(1677) <= "0000000000000000";
ram(1678) <= "0000000000000000";
ram(1679) <= "0000000000000000";
ram(1680) <= "0000000000000000";
ram(1681) <= "0000000000000000";
ram(1682) <= "0000000000000000";
ram(1683) <= "0000000000000000";
ram(1684) <= "0000000000000000";
ram(1685) <= "0000000000000000";
ram(1686) <= "0000000000000000";
ram(1687) <= "0000000000000000";
ram(1688) <= "0000000000000000";
ram(1689) <= "0000000000000000";
ram(1690) <= "0000000000000000";
ram(1691) <= "0000000000000000";
ram(1692) <= "0000000000000000";
ram(1693) <= "0000000000000000";
ram(1694) <= "0000000000000000";
ram(1695) <= "0000000000000000";
ram(1696) <= "0000000000000000";
ram(1697) <= "0000000000000000";
ram(1698) <= "0000000000000000";
ram(1699) <= "0000000000000000";
ram(1700) <= "0000000000000000";
ram(1701) <= "0000000000000000";
ram(1702) <= "0000000000000000";
ram(1703) <= "0000000000000000";
ram(1704) <= "0000000000000000";
ram(1705) <= "0000000000000000";
ram(1706) <= "0000000000000000";
ram(1707) <= "0000000000000000";
ram(1708) <= "0000000000000000";
ram(1709) <= "0000000000000000";
ram(1710) <= "0000000000000000";
ram(1711) <= "0000000000000000";
ram(1712) <= "0000000000000000";
ram(1713) <= "0000000000000000";
ram(1714) <= "0000000000000000";
ram(1715) <= "0000000000000000";
ram(1716) <= "0000000000000000";
ram(1717) <= "0000000000000000";
ram(1718) <= "0000000000000000";
ram(1719) <= "0000000000000000";
ram(1720) <= "0000000000000000";
ram(1721) <= "0000000000000000";
ram(1722) <= "0000000000000000";
ram(1723) <= "0000000000000000";
ram(1724) <= "0000000000000000";
ram(1725) <= "0000000000000000";
ram(1726) <= "0000000000000000";
ram(1727) <= "0000000000000000";
ram(1728) <= "0000000000000000";
ram(1729) <= "0000000000000000";
ram(1730) <= "0000000000000000";
ram(1731) <= "0000000000000000";
ram(1732) <= "0000000000000000";
ram(1733) <= "0000000000000000";
ram(1734) <= "0000000000000000";
ram(1735) <= "0000000000000000";
ram(1736) <= "0000000000000000";
ram(1737) <= "0000000000000000";
ram(1738) <= "0000000000000000";
ram(1739) <= "0000000000000000";
ram(1740) <= "0000000000000000";
ram(1741) <= "0000000000000000";
ram(1742) <= "0000000000000000";
ram(1743) <= "0000000000000000";
ram(1744) <= "0000000000000000";
ram(1745) <= "0000000000000000";
ram(1746) <= "0000000000000000";
ram(1747) <= "0000000000000000";
ram(1748) <= "0000000000000000";
ram(1749) <= "0000000000000000";
ram(1750) <= "0000000000000000";
ram(1751) <= "0000000000000000";
ram(1752) <= "0000000000000000";
ram(1753) <= "0000000000000000";
ram(1754) <= "0000000000000000";
ram(1755) <= "0000000000000000";
ram(1756) <= "0000000000000000";
ram(1757) <= "0000000000000000";
ram(1758) <= "0000000000000000";
ram(1759) <= "0000000000000000";
ram(1760) <= "0000000000000000";
ram(1761) <= "0000000000000000";
ram(1762) <= "0000000000000000";
ram(1763) <= "0000000000000000";
ram(1764) <= "0000000000000000";
ram(1765) <= "0000000000000000";
ram(1766) <= "0000000000000000";
ram(1767) <= "0000000000000000";
ram(1768) <= "0000000000000000";
ram(1769) <= "0000000000000000";
ram(1770) <= "0000000000000000";
ram(1771) <= "0000000000000000";
ram(1772) <= "0000000000000000";
ram(1773) <= "0000000000000000";
ram(1774) <= "0000000000000000";
ram(1775) <= "0000000000000000";
ram(1776) <= "0000000000000000";
ram(1777) <= "0000000000000000";
ram(1778) <= "0000000000000000";
ram(1779) <= "0000000000000000";
ram(1780) <= "0000000000000000";
ram(1781) <= "0000000000000000";
ram(1782) <= "0000000000000000";
ram(1783) <= "0000000000000000";
ram(1784) <= "0000000000000000";
ram(1785) <= "0000000000000000";
ram(1786) <= "0000000000000000";
ram(1787) <= "0000000000000000";
ram(1788) <= "0000000000000000";
ram(1789) <= "0000000000000000";
ram(1790) <= "0000000000000000";
ram(1791) <= "0000000000000000";
ram(1792) <= "0000000000000000";
ram(1793) <= "0000000000000000";
ram(1794) <= "0000000000000000";
ram(1795) <= "0000000000000000";
ram(1796) <= "0000000000000000";
ram(1797) <= "0000000000000000";
ram(1798) <= "0000000000000000";
ram(1799) <= "0000000000000000";
ram(1800) <= "0000000000000000";
ram(1801) <= "0000000000000000";
ram(1802) <= "0000000000000000";
ram(1803) <= "0000000000000000";
ram(1804) <= "0000000000000000";
ram(1805) <= "0000000000000000";
ram(1806) <= "0000000000000000";
ram(1807) <= "0000000000000000";
ram(1808) <= "0000000000000000";
ram(1809) <= "0000000000000000";
ram(1810) <= "0000000000000000";
ram(1811) <= "0000000000000000";
ram(1812) <= "0000000000000000";
ram(1813) <= "0000000000000000";
ram(1814) <= "0000000000000000";
ram(1815) <= "0000000000000000";
ram(1816) <= "0000000000000000";
ram(1817) <= "0000000000000000";
ram(1818) <= "0000000000000000";
ram(1819) <= "0000000000000000";
ram(1820) <= "0000000000000000";
ram(1821) <= "0000000000000000";
ram(1822) <= "0000000000000000";
ram(1823) <= "0000000000000000";
ram(1824) <= "0000000000000000";
ram(1825) <= "0000000000000000";
ram(1826) <= "0000000000000000";
ram(1827) <= "0000000000000000";
ram(1828) <= "0000000000000000";
ram(1829) <= "0000000000000000";
ram(1830) <= "0000000000000000";
ram(1831) <= "0000000000000000";
ram(1832) <= "0000000000000000";
ram(1833) <= "0000000000000000";
ram(1834) <= "0000000000000000";
ram(1835) <= "0000000000000000";
ram(1836) <= "0000000000000000";
ram(1837) <= "0000000000000000";
ram(1838) <= "0000000000000000";
ram(1839) <= "0000000000000000";
ram(1840) <= "0000000000000000";
ram(1841) <= "0000000000000000";
ram(1842) <= "0000000000000000";
ram(1843) <= "0000000000000000";
ram(1844) <= "0000000000000000";
ram(1845) <= "0000000000000000";
ram(1846) <= "0000000000000000";
ram(1847) <= "0000000000000000";
ram(1848) <= "0000000000000000";
ram(1849) <= "0000000000000000";
ram(1850) <= "0000000000000000";
ram(1851) <= "0000000000000000";
ram(1852) <= "0000000000000000";
ram(1853) <= "0000000000000000";
ram(1854) <= "0000000000000000";
ram(1855) <= "0000000000000000";
ram(1856) <= "0000000000000000";
ram(1857) <= "0000000000000000";
ram(1858) <= "0000000000000000";
ram(1859) <= "0000000000000000";
ram(1860) <= "0000000000000000";
ram(1861) <= "0000000000000000";
ram(1862) <= "0000000000000000";
ram(1863) <= "0000000000000000";
ram(1864) <= "0000000000000000";
ram(1865) <= "0000000000000000";
ram(1866) <= "0000000000000000";
ram(1867) <= "0000000000000000";
ram(1868) <= "0000000000000000";
ram(1869) <= "0000000000000000";
ram(1870) <= "0000000000000000";
ram(1871) <= "0000000000000000";
ram(1872) <= "0000000000000000";
ram(1873) <= "0000000000000000";
ram(1874) <= "0000000000000000";
ram(1875) <= "0000000000000000";
ram(1876) <= "0000000000000000";
ram(1877) <= "0000000000000000";
ram(1878) <= "0000000000000000";
ram(1879) <= "0000000000000000";
ram(1880) <= "0000000000000000";
ram(1881) <= "0000000000000000";
ram(1882) <= "0000000000000000";
ram(1883) <= "0000000000000000";
ram(1884) <= "0000000000000000";
ram(1885) <= "0000000000000000";
ram(1886) <= "0000000000000000";
ram(1887) <= "0000000000000000";
ram(1888) <= "0000000000000000";
ram(1889) <= "0000000000000000";
ram(1890) <= "0000000000000000";
ram(1891) <= "0000000000000000";
ram(1892) <= "0000000000000000";
ram(1893) <= "0000000000000000";
ram(1894) <= "0000000000000000";
ram(1895) <= "0000000000000000";
ram(1896) <= "0000000000000000";
ram(1897) <= "0000000000000000";
ram(1898) <= "0000000000000000";
ram(1899) <= "0000000000000000";
ram(1900) <= "0000000000000000";
ram(1901) <= "0000000000000000";
ram(1902) <= "0000000000000000";
ram(1903) <= "0000000000000000";
ram(1904) <= "0000000000000000";
ram(1905) <= "0000000000000000";
ram(1906) <= "0000000000000000";
ram(1907) <= "0000000000000000";
ram(1908) <= "0000000000000000";
ram(1909) <= "0000000000000000";
ram(1910) <= "0000000000000000";
ram(1911) <= "0000000000000000";
ram(1912) <= "0000000000000000";
ram(1913) <= "0000000000000000";
ram(1914) <= "0000000000000000";
ram(1915) <= "0000000000000000";
ram(1916) <= "0000000000000000";
ram(1917) <= "0000000000000000";
ram(1918) <= "0000000000000000";
ram(1919) <= "0000000000000000";
ram(1920) <= "0000000000000000";
ram(1921) <= "0000000000000000";
ram(1922) <= "0000000000000000";
ram(1923) <= "0000000000000000";
ram(1924) <= "0000000000000000";
ram(1925) <= "0000000000000000";
ram(1926) <= "0000000000000000";
ram(1927) <= "0000000000000000";
ram(1928) <= "0000000000000000";
ram(1929) <= "0000000000000000";
ram(1930) <= "0000000000000000";
ram(1931) <= "0000000000000000";
ram(1932) <= "0000000000000000";
ram(1933) <= "0000000000000000";
ram(1934) <= "0000000000000000";
ram(1935) <= "0000000000000000";
ram(1936) <= "0000000000000000";
ram(1937) <= "0000000000000000";
ram(1938) <= "0000000000000000";
ram(1939) <= "0000000000000000";
ram(1940) <= "0000000000000000";
ram(1941) <= "0000000000000000";
ram(1942) <= "0000000000000000";
ram(1943) <= "0000000000000000";
ram(1944) <= "0000000000000000";
ram(1945) <= "0000000000000000";
ram(1946) <= "0000000000000000";
ram(1947) <= "0000000000000000";
ram(1948) <= "0000000000000000";
ram(1949) <= "0000000000000000";
ram(1950) <= "0000000000000000";
ram(1951) <= "0000000000000000";
ram(1952) <= "0000000000000000";
ram(1953) <= "0000000000000000";
ram(1954) <= "0000000000000000";
ram(1955) <= "0000000000000000";
ram(1956) <= "0000000000000000";
ram(1957) <= "0000000000000000";
ram(1958) <= "0000000000000000";
ram(1959) <= "0000000000000000";
ram(1960) <= "0000000000000000";
ram(1961) <= "0000000000000000";
ram(1962) <= "0000000000000000";
ram(1963) <= "0000000000000000";
ram(1964) <= "0000000000000000";
ram(1965) <= "0000000000000000";
ram(1966) <= "0000000000000000";
ram(1967) <= "0000000000000000";
ram(1968) <= "0000000000000000";
ram(1969) <= "0000000000000000";
ram(1970) <= "0000000000000000";
ram(1971) <= "0000000000000000";
ram(1972) <= "0000000000000000";
ram(1973) <= "0000000000000000";
ram(1974) <= "0000000000000000";
ram(1975) <= "0000000000000000";
ram(1976) <= "0000000000000000";
ram(1977) <= "0000000000000000";
ram(1978) <= "0000000000000000";
ram(1979) <= "0000000000000000";
ram(1980) <= "0000000000000000";
ram(1981) <= "0000000000000000";
ram(1982) <= "0000000000000000";
ram(1983) <= "0000000000000000";
ram(1984) <= "0000000000000000";
ram(1985) <= "0000000000000000";
ram(1986) <= "0000000000000000";
ram(1987) <= "0000000000000000";
ram(1988) <= "0000000000000000";
ram(1989) <= "0000000000000000";
ram(1990) <= "0000000000000000";
ram(1991) <= "0000000000000000";
ram(1992) <= "0000000000000000";
ram(1993) <= "0000000000000000";
ram(1994) <= "0000000000000000";
ram(1995) <= "0000000000000000";
ram(1996) <= "0000000000000000";
ram(1997) <= "0000000000000000";
ram(1998) <= "0000000000000000";
ram(1999) <= "0000000000000000";
ram(2000) <= "0000000000000000";
ram(2001) <= "0000000000000000";
ram(2002) <= "0000000000000000";
ram(2003) <= "0000000000000000";
ram(2004) <= "0000000000000000";
ram(2005) <= "0000000000000000";
ram(2006) <= "0000000000000000";
ram(2007) <= "0000000000000000";
ram(2008) <= "0000000000000000";
ram(2009) <= "0000000000000000";
ram(2010) <= "0000000000000000";
ram(2011) <= "0000000000000000";
ram(2012) <= "0000000000000000";
ram(2013) <= "0000000000000000";
ram(2014) <= "0000000000000000";
ram(2015) <= "0000000000000000";
ram(2016) <= "0000000000000000";
ram(2017) <= "0000000000000000";
ram(2018) <= "0000000000000000";
ram(2019) <= "0000000000000000";
ram(2020) <= "0000000000000000";
ram(2021) <= "0000000000000000";
ram(2022) <= "0000000000000000";
ram(2023) <= "0000000000000000";
ram(2024) <= "0000000000000000";
ram(2025) <= "0000000000000000";
ram(2026) <= "0000000000000000";
ram(2027) <= "0000000000000000";
ram(2028) <= "0000000000000000";
ram(2029) <= "0000000000000000";
ram(2030) <= "0000000000000000";
ram(2031) <= "0000000000000000";
ram(2032) <= "0000000000000000";
ram(2033) <= "0000000000000000";
ram(2034) <= "0000000000000000";
ram(2035) <= "0000000000000000";
ram(2036) <= "0000000000000000";
ram(2037) <= "0000000000000000";
ram(2038) <= "0000000000000000";
ram(2039) <= "0000000000000000";
ram(2040) <= "0000000000000000";
ram(2041) <= "0000000000000000";
ram(2042) <= "0000000000000000";
ram(2043) <= "0000000000000000";
ram(2044) <= "0000000000000000";
ram(2045) <= "0000000000000000";
ram(2046) <= "0000000000000000";
ram(2047) <= "0000000000000000";
ram(2048) <= "0000000000000000";
ram(2049) <= "0000000000000000";
ram(2050) <= "0000000000000000";
ram(2051) <= "0000000000000000";
ram(2052) <= "0000000000000000";
ram(2053) <= "0000000000000000";
ram(2054) <= "0000000000000000";
ram(2055) <= "0000000000000000";
ram(2056) <= "0000000000000000";
ram(2057) <= "0000000000000000";
ram(2058) <= "0000000000000000";
ram(2059) <= "0000000000000000";
ram(2060) <= "0000000000000000";
ram(2061) <= "0000000000000000";
ram(2062) <= "0000000000000000";
ram(2063) <= "0000000000000000";
ram(2064) <= "0000000000000000";
ram(2065) <= "0000000000000000";
ram(2066) <= "0000000000000000";
ram(2067) <= "0000000000000000";
ram(2068) <= "0000000000000000";
ram(2069) <= "0000000000000000";
ram(2070) <= "0000000000000000";
ram(2071) <= "0000000000000000";
ram(2072) <= "0000000000000000";
ram(2073) <= "0000000000000000";
ram(2074) <= "0000000000000000";
ram(2075) <= "0000000000000000";
ram(2076) <= "0000000000000000";
ram(2077) <= "0000000000000000";
ram(2078) <= "0000000000000000";
ram(2079) <= "0000000000000000";
ram(2080) <= "0000000000000000";
ram(2081) <= "0000000000000000";
ram(2082) <= "0000000000000000";
ram(2083) <= "0000000000000000";
ram(2084) <= "0000000000000000";
ram(2085) <= "0000000000000000";
ram(2086) <= "0000000000000000";
ram(2087) <= "0000000000000000";
ram(2088) <= "0000000000000000";
ram(2089) <= "0000000000000000";
ram(2090) <= "0000000000000000";
ram(2091) <= "0000000000000000";
ram(2092) <= "0000000000000000";
ram(2093) <= "0000000000000000";
ram(2094) <= "0000000000000000";
ram(2095) <= "0000000000000000";
ram(2096) <= "0000000000000000";
ram(2097) <= "0000000000000000";
ram(2098) <= "0000000000000000";
ram(2099) <= "0000000000000000";
ram(2100) <= "0000000000000000";
ram(2101) <= "0000000000000000";
ram(2102) <= "0000000000000000";
ram(2103) <= "0000000000000000";
ram(2104) <= "0000000000000000";
ram(2105) <= "0000000000000000";
ram(2106) <= "0000000000000000";
ram(2107) <= "0000000000000000";
ram(2108) <= "0000000000000000";
ram(2109) <= "0000000000000000";
ram(2110) <= "0000000000000000";
ram(2111) <= "0000000000000000";
ram(2112) <= "0000000000000000";
ram(2113) <= "0000000000000000";
ram(2114) <= "0000000000000000";
ram(2115) <= "0000000000000000";
ram(2116) <= "0000000000000000";
ram(2117) <= "0000000000000000";
ram(2118) <= "0000000000000000";
ram(2119) <= "0000000000000000";
ram(2120) <= "0000000000000000";
ram(2121) <= "0000000000000000";
ram(2122) <= "0000000000000000";
ram(2123) <= "0000000000000000";
ram(2124) <= "0000000000000000";
ram(2125) <= "0000000000000000";
ram(2126) <= "0000000000000000";
ram(2127) <= "0000000000000000";
ram(2128) <= "0000000000000000";
ram(2129) <= "0000000000000000";
ram(2130) <= "0000000000000000";
ram(2131) <= "0000000000000000";
ram(2132) <= "0000000000000000";
ram(2133) <= "0000000000000000";
ram(2134) <= "0000000000000000";
ram(2135) <= "0000000000000000";
ram(2136) <= "0000000000000000";
ram(2137) <= "0000000000000000";
ram(2138) <= "0000000000000000";
ram(2139) <= "0000000000000000";
ram(2140) <= "0000000000000000";
ram(2141) <= "0000000000000000";
ram(2142) <= "0000000000000000";
ram(2143) <= "0000000000000000";
ram(2144) <= "0000000000000000";
ram(2145) <= "0000000000000000";
ram(2146) <= "0000000000000000";
ram(2147) <= "0000000000000000";
ram(2148) <= "0000000000000000";
ram(2149) <= "0000000000000000";
ram(2150) <= "0000000000000000";
ram(2151) <= "0000000000000000";
ram(2152) <= "0000000000000000";
ram(2153) <= "0000000000000000";
ram(2154) <= "0000000000000000";
ram(2155) <= "0000000000000000";
ram(2156) <= "0000000000000000";
ram(2157) <= "0000000000000000";
ram(2158) <= "0000000000000000";
ram(2159) <= "0000000000000000";
ram(2160) <= "0000000000000000";
ram(2161) <= "0000000000000000";
ram(2162) <= "0000000000000000";
ram(2163) <= "0000000000000000";
ram(2164) <= "0000000000000000";
ram(2165) <= "0000000000000000";
ram(2166) <= "0000000000000000";
ram(2167) <= "0000000000000000";
ram(2168) <= "0000000000000000";
ram(2169) <= "0000000000000000";
ram(2170) <= "0000000000000000";
ram(2171) <= "0000000000000000";
ram(2172) <= "0000000000000000";
ram(2173) <= "0000000000000000";
ram(2174) <= "0000000000000000";
ram(2175) <= "0000000000000000";
ram(2176) <= "0000000000000000";
ram(2177) <= "0000000000000000";
ram(2178) <= "0000000000000000";
ram(2179) <= "0000000000000000";
ram(2180) <= "0000000000000000";
ram(2181) <= "0000000000000000";
ram(2182) <= "0000000000000000";
ram(2183) <= "0000000000000000";
ram(2184) <= "0000000000000000";
ram(2185) <= "0000000000000000";
ram(2186) <= "0000000000000000";
ram(2187) <= "0000000000000000";
ram(2188) <= "0000000000000000";
ram(2189) <= "0000000000000000";
ram(2190) <= "0000000000000000";
ram(2191) <= "0000000000000000";
ram(2192) <= "0000000000000000";
ram(2193) <= "0000000000000000";
ram(2194) <= "0000000000000000";
ram(2195) <= "0000000000000000";
ram(2196) <= "0000000000000000";
ram(2197) <= "0000000000000000";
ram(2198) <= "0000000000000000";
ram(2199) <= "0000000000000000";
ram(2200) <= "0000000000000000";
ram(2201) <= "0000000000000000";
ram(2202) <= "0000000000000000";
ram(2203) <= "0000000000000000";
ram(2204) <= "0000000000000000";
ram(2205) <= "0000000000000000";
ram(2206) <= "0000000000000000";
ram(2207) <= "0000000000000000";
ram(2208) <= "0000000000000000";
ram(2209) <= "0000000000000000";
ram(2210) <= "0000000000000000";
ram(2211) <= "0000000000000000";
ram(2212) <= "0000000000000000";
ram(2213) <= "0000000000000000";
ram(2214) <= "0000000000000000";
ram(2215) <= "0000000000000000";
ram(2216) <= "0000000000000000";
ram(2217) <= "0000000000000000";
ram(2218) <= "0000000000000000";
ram(2219) <= "0000000000000000";
ram(2220) <= "0000000000000000";
ram(2221) <= "0000000000000000";
ram(2222) <= "0000000000000000";
ram(2223) <= "0000000000000000";
ram(2224) <= "0000000000000000";
ram(2225) <= "0000000000000000";
ram(2226) <= "0000000000000000";
ram(2227) <= "0000000000000000";
ram(2228) <= "0000000000000000";
ram(2229) <= "0000000000000000";
ram(2230) <= "0000000000000000";
ram(2231) <= "0000000000000000";
ram(2232) <= "0000000000000000";
ram(2233) <= "0000000000000000";
ram(2234) <= "0000000000000000";
ram(2235) <= "0000000000000000";
ram(2236) <= "0000000000000000";
ram(2237) <= "0000000000000000";
ram(2238) <= "0000000000000000";
ram(2239) <= "0000000000000000";
ram(2240) <= "0000000000000000";
ram(2241) <= "0000000000000000";
ram(2242) <= "0000000000000000";
ram(2243) <= "0000000000000000";
ram(2244) <= "0000000000000000";
ram(2245) <= "0000000000000000";
ram(2246) <= "0000000000000000";
ram(2247) <= "0000000000000000";
ram(2248) <= "0000000000000000";
ram(2249) <= "0000000000000000";
ram(2250) <= "0000000000000000";
ram(2251) <= "0000000000000000";
ram(2252) <= "0000000000000000";
ram(2253) <= "0000000000000000";
ram(2254) <= "0000000000000000";
ram(2255) <= "0000000000000000";
ram(2256) <= "0000000000000000";
ram(2257) <= "0000000000000000";
ram(2258) <= "0000000000000000";
ram(2259) <= "0000000000000000";
ram(2260) <= "0000000000000000";
ram(2261) <= "0000000000000000";
ram(2262) <= "0000000000000000";
ram(2263) <= "0000000000000000";
ram(2264) <= "0000000000000000";
ram(2265) <= "0000000000000000";
ram(2266) <= "0000000000000000";
ram(2267) <= "0000000000000000";
ram(2268) <= "0000000000000000";
ram(2269) <= "0000000000000000";
ram(2270) <= "0000000000000000";
ram(2271) <= "0000000000000000";
ram(2272) <= "0000000000000000";
ram(2273) <= "0000000000000000";
ram(2274) <= "0000000000000000";
ram(2275) <= "0000000000000000";
ram(2276) <= "0000000000000000";
ram(2277) <= "0000000000000000";
ram(2278) <= "0000000000000000";
ram(2279) <= "0000000000000000";
ram(2280) <= "0000000000000000";
ram(2281) <= "0000000000000000";
ram(2282) <= "0000000000000000";
ram(2283) <= "0000000000000000";
ram(2284) <= "0000000000000000";
ram(2285) <= "0000000000000000";
ram(2286) <= "0000000000000000";
ram(2287) <= "0000000000000000";
ram(2288) <= "0000000000000000";
ram(2289) <= "0000000000000000";
ram(2290) <= "0000000000000000";
ram(2291) <= "0000000000000000";
ram(2292) <= "0000000000000000";
ram(2293) <= "0000000000000000";
ram(2294) <= "0000000000000000";
ram(2295) <= "0000000000000000";
ram(2296) <= "0000000000000000";
ram(2297) <= "0000000000000000";
ram(2298) <= "0000000000000000";
ram(2299) <= "0000000000000000";
ram(2300) <= "0000000000000000";
ram(2301) <= "0000000000000000";
ram(2302) <= "0000000000000000";
ram(2303) <= "0000000000000000";
ram(2304) <= "0000000000000000";
ram(2305) <= "0000000000000000";
ram(2306) <= "0000000000000000";
ram(2307) <= "0000000000000000";
ram(2308) <= "0000000000000000";
ram(2309) <= "0000000000000000";
ram(2310) <= "0000000000000000";
ram(2311) <= "0000000000000000";
ram(2312) <= "0000000000000000";
ram(2313) <= "0000000000000000";
ram(2314) <= "0000000000000000";
ram(2315) <= "0000000000000000";
ram(2316) <= "0000000000000000";
ram(2317) <= "0000000000000000";
ram(2318) <= "0000000000000000";
ram(2319) <= "0000000000000000";
ram(2320) <= "0000000000000000";
ram(2321) <= "0000000000000000";
ram(2322) <= "0000000000000000";
ram(2323) <= "0000000000000000";
ram(2324) <= "0000000000000000";
ram(2325) <= "0000000000000000";
ram(2326) <= "0000000000000000";
ram(2327) <= "0000000000000000";
ram(2328) <= "0000000000000000";
ram(2329) <= "0000000000000000";
ram(2330) <= "0000000000000000";
ram(2331) <= "0000000000000000";
ram(2332) <= "0000000000000000";
ram(2333) <= "0000000000000000";
ram(2334) <= "0000000000000000";
ram(2335) <= "0000000000000000";
ram(2336) <= "0000000000000000";
ram(2337) <= "0000000000000000";
ram(2338) <= "0000000000000000";
ram(2339) <= "0000000000000000";
ram(2340) <= "0000000000000000";
ram(2341) <= "0000000000000000";
ram(2342) <= "0000000000000000";
ram(2343) <= "0000000000000000";
ram(2344) <= "0000000000000000";
ram(2345) <= "0000000000000000";
ram(2346) <= "0000000000000000";
ram(2347) <= "0000000000000000";
ram(2348) <= "0000000000000000";
ram(2349) <= "0000000000000000";
ram(2350) <= "0000000000000000";
ram(2351) <= "0000000000000000";
ram(2352) <= "0000000000000000";
ram(2353) <= "0000000000000000";
ram(2354) <= "0000000000000000";
ram(2355) <= "0000000000000000";
ram(2356) <= "0000000000000000";
ram(2357) <= "0000000000000000";
ram(2358) <= "0000000000000000";
ram(2359) <= "0000000000000000";
ram(2360) <= "0000000000000000";
ram(2361) <= "0000000000000000";
ram(2362) <= "0000000000000000";
ram(2363) <= "0000000000000000";
ram(2364) <= "0000000000000000";
ram(2365) <= "0000000000000000";
ram(2366) <= "0000000000000000";
ram(2367) <= "0000000000000000";
ram(2368) <= "0000000000000000";
ram(2369) <= "0000000000000000";
ram(2370) <= "0000000000000000";
ram(2371) <= "0000000000000000";
ram(2372) <= "0000000000000000";
ram(2373) <= "0000000000000000";
ram(2374) <= "0000000000000000";
ram(2375) <= "0000000000000000";
ram(2376) <= "0000000000000000";
ram(2377) <= "0000000000000000";
ram(2378) <= "0000000000000000";
ram(2379) <= "0000000000000000";
ram(2380) <= "0000000000000000";
ram(2381) <= "0000000000000000";
ram(2382) <= "0000000000000000";
ram(2383) <= "0000000000000000";
ram(2384) <= "0000000000000000";
ram(2385) <= "0000000000000000";
ram(2386) <= "0000000000000000";
ram(2387) <= "0000000000000000";
ram(2388) <= "0000000000000000";
ram(2389) <= "0000000000000000";
ram(2390) <= "0000000000000000";
ram(2391) <= "0000000000000000";
ram(2392) <= "0000000000000000";
ram(2393) <= "0000000000000000";
ram(2394) <= "0000000000000000";
ram(2395) <= "0000000000000000";
ram(2396) <= "0000000000000000";
ram(2397) <= "0000000000000000";
ram(2398) <= "0000000000000000";
ram(2399) <= "0000000000000000";
ram(2400) <= "0000000000000000";
ram(2401) <= "0000000000000000";
ram(2402) <= "0000000000000000";
ram(2403) <= "0000000000000000";
ram(2404) <= "0000000000000000";
ram(2405) <= "0000000000000000";
ram(2406) <= "0000000000000000";
ram(2407) <= "0000000000000000";
ram(2408) <= "0000000000000000";
ram(2409) <= "0000000000000000";
ram(2410) <= "0000000000000000";
ram(2411) <= "0000000000000000";
ram(2412) <= "0000000000000000";
ram(2413) <= "0000000000000000";
ram(2414) <= "0000000000000000";
ram(2415) <= "0000000000000000";
ram(2416) <= "0000000000000000";
ram(2417) <= "0000000000000000";
ram(2418) <= "0000000000000000";
ram(2419) <= "0000000000000000";
ram(2420) <= "0000000000000000";
ram(2421) <= "0000000000000000";
ram(2422) <= "0000000000000000";
ram(2423) <= "0000000000000000";
ram(2424) <= "0000000000000000";
ram(2425) <= "0000000000000000";
ram(2426) <= "0000000000000000";
ram(2427) <= "0000000000000000";
ram(2428) <= "0000000000000000";
ram(2429) <= "0000000000000000";
ram(2430) <= "0000000000000000";
ram(2431) <= "0000000000000000";
ram(2432) <= "0000000000000000";
ram(2433) <= "0000000000000000";
ram(2434) <= "0000000000000000";
ram(2435) <= "0000000000000000";
ram(2436) <= "0000000000000000";
ram(2437) <= "0000000000000000";
ram(2438) <= "0000000000000000";
ram(2439) <= "0000000000000000";
ram(2440) <= "0000000000000000";
ram(2441) <= "0000000000000000";
ram(2442) <= "0000000000000000";
ram(2443) <= "0000000000000000";
ram(2444) <= "0000000000000000";
ram(2445) <= "0000000000000000";
ram(2446) <= "0000000000000000";
ram(2447) <= "0000000000000000";
ram(2448) <= "0000000000000000";
ram(2449) <= "0000000000000000";
ram(2450) <= "0000000000000000";
ram(2451) <= "0000000000000000";
ram(2452) <= "0000000000000000";
ram(2453) <= "0000000000000000";
ram(2454) <= "0000000000000000";
ram(2455) <= "0000000000000000";
ram(2456) <= "0000000000000000";
ram(2457) <= "0000000000000000";
ram(2458) <= "0000000000000000";
ram(2459) <= "0000000000000000";
ram(2460) <= "0000000000000000";
ram(2461) <= "0000000000000000";
ram(2462) <= "0000000000000000";
ram(2463) <= "0000000000000000";
ram(2464) <= "0000000000000000";
ram(2465) <= "0000000000000000";
ram(2466) <= "0000000000000000";
ram(2467) <= "0000000000000000";
ram(2468) <= "0000000000000000";
ram(2469) <= "0000000000000000";
ram(2470) <= "0000000000000000";
ram(2471) <= "0000000000000000";
ram(2472) <= "0000000000000000";
ram(2473) <= "0000000000000000";
ram(2474) <= "0000000000000000";
ram(2475) <= "0000000000000000";
ram(2476) <= "0000000000000000";
ram(2477) <= "0000000000000000";
ram(2478) <= "0000000000000000";
ram(2479) <= "0000000000000000";
ram(2480) <= "0000000000000000";
ram(2481) <= "0000000000000000";
ram(2482) <= "0000000000000000";
ram(2483) <= "0000000000000000";
ram(2484) <= "0000000000000000";
ram(2485) <= "0000000000000000";
ram(2486) <= "0000000000000000";
ram(2487) <= "0000000000000000";
ram(2488) <= "0000000000000000";
ram(2489) <= "0000000000000000";
ram(2490) <= "0000000000000000";
ram(2491) <= "0000000000000000";
ram(2492) <= "0000000000000000";
ram(2493) <= "0000000000000000";
ram(2494) <= "0000000000000000";
ram(2495) <= "0000000000000000";
ram(2496) <= "0000000000000000";
ram(2497) <= "0000000000000000";
ram(2498) <= "0000000000000000";
ram(2499) <= "0000000000000000";
ram(2500) <= "0000000000000000";
ram(2501) <= "0000000000000000";
ram(2502) <= "0000000000000000";
ram(2503) <= "0000000000000000";
ram(2504) <= "0000000000000000";
ram(2505) <= "0000000000000000";
ram(2506) <= "0000000000000000";
ram(2507) <= "0000000000000000";
ram(2508) <= "0000000000000000";
ram(2509) <= "0000000000000000";
ram(2510) <= "0000000000000000";
ram(2511) <= "0000000000000000";
ram(2512) <= "0000000000000000";
ram(2513) <= "0000000000000000";
ram(2514) <= "0000000000000000";
ram(2515) <= "0000000000000000";
ram(2516) <= "0000000000000000";
ram(2517) <= "0000000000000000";
ram(2518) <= "0000000000000000";
ram(2519) <= "0000000000000000";
ram(2520) <= "0000000000000000";
ram(2521) <= "0000000000000000";
ram(2522) <= "0000000000000000";
ram(2523) <= "0000000000000000";
ram(2524) <= "0000000000000000";
ram(2525) <= "0000000000000000";
ram(2526) <= "0000000000000000";
ram(2527) <= "0000000000000000";
ram(2528) <= "0000000000000000";
ram(2529) <= "0000000000000000";
ram(2530) <= "0000000000000000";
ram(2531) <= "0000000000000000";
ram(2532) <= "0000000000000000";
ram(2533) <= "0000000000000000";
ram(2534) <= "0000000000000000";
ram(2535) <= "0000000000000000";
ram(2536) <= "0000000000000000";
ram(2537) <= "0000000000000000";
ram(2538) <= "0000000000000000";
ram(2539) <= "0000000000000000";
ram(2540) <= "0000000000000000";
ram(2541) <= "0000000000000000";
ram(2542) <= "0000000000000000";
ram(2543) <= "0000000000000000";
ram(2544) <= "0000000000000000";
ram(2545) <= "0000000000000000";
ram(2546) <= "0000000000000000";
ram(2547) <= "0000000000000000";
ram(2548) <= "0000000000000000";
ram(2549) <= "0000000000000000";
ram(2550) <= "0000000000000000";
ram(2551) <= "0000000000000000";
ram(2552) <= "0000000000000000";
ram(2553) <= "0000000000000000";
ram(2554) <= "0000000000000000";
ram(2555) <= "0000000000000000";
ram(2556) <= "0000000000000000";
ram(2557) <= "0000000000000000";
ram(2558) <= "0000000000000000";
ram(2559) <= "0000000000000000";
ram(2560) <= "0000000000000000";
ram(2561) <= "0000000000000000";
ram(2562) <= "0000000000000000";
ram(2563) <= "0000000000000000";
ram(2564) <= "0000000000000000";
ram(2565) <= "0000000000000000";
ram(2566) <= "0000000000000000";
ram(2567) <= "0000000000000000";
ram(2568) <= "0000000000000000";
ram(2569) <= "0000000000000000";
ram(2570) <= "0000000000000000";
ram(2571) <= "0000000000000000";
ram(2572) <= "0000000000000000";
ram(2573) <= "0000000000000000";
ram(2574) <= "0000000000000000";
ram(2575) <= "0000000000000000";
ram(2576) <= "0000000000000000";
ram(2577) <= "0000000000000000";
ram(2578) <= "0000000000000000";
ram(2579) <= "0000000000000000";
ram(2580) <= "0000000000000000";
ram(2581) <= "0000000000000000";
ram(2582) <= "0000000000000000";
ram(2583) <= "0000000000000000";
ram(2584) <= "0000000000000000";
ram(2585) <= "0000000000000000";
ram(2586) <= "0000000000000000";
ram(2587) <= "0000000000000000";
ram(2588) <= "0000000000000000";
ram(2589) <= "0000000000000000";
ram(2590) <= "0000000000000000";
ram(2591) <= "0000000000000000";
ram(2592) <= "0000000000000000";
ram(2593) <= "0000000000000000";
ram(2594) <= "0000000000000000";
ram(2595) <= "0000000000000000";
ram(2596) <= "0000000000000000";
ram(2597) <= "0000000000000000";
ram(2598) <= "0000000000000000";
ram(2599) <= "0000000000000000";
ram(2600) <= "0000000000000000";
ram(2601) <= "0000000000000000";
ram(2602) <= "0000000000000000";
ram(2603) <= "0000000000000000";
ram(2604) <= "0000000000000000";
ram(2605) <= "0000000000000000";
ram(2606) <= "0000000000000000";
ram(2607) <= "0000000000000000";
ram(2608) <= "0000000000000000";
ram(2609) <= "0000000000000000";
ram(2610) <= "0000000000000000";
ram(2611) <= "0000000000000000";
ram(2612) <= "0000000000000000";
ram(2613) <= "0000000000000000";
ram(2614) <= "0000000000000000";
ram(2615) <= "0000000000000000";
ram(2616) <= "0000000000000000";
ram(2617) <= "0000000000000000";
ram(2618) <= "0000000000000000";
ram(2619) <= "0000000000000000";
ram(2620) <= "0000000000000000";
ram(2621) <= "0000000000000000";
ram(2622) <= "0000000000000000";
ram(2623) <= "0000000000000000";
ram(2624) <= "0000000000000000";
ram(2625) <= "0000000000000000";
ram(2626) <= "0000000000000000";
ram(2627) <= "0000000000000000";
ram(2628) <= "0000000000000000";
ram(2629) <= "0000000000000000";
ram(2630) <= "0000000000000000";
ram(2631) <= "0000000000000000";
ram(2632) <= "0000000000000000";
ram(2633) <= "0000000000000000";
ram(2634) <= "0000000000000000";
ram(2635) <= "0000000000000000";
ram(2636) <= "0000000000000000";
ram(2637) <= "0000000000000000";
ram(2638) <= "0000000000000000";
ram(2639) <= "0000000000000000";
ram(2640) <= "0000000000000000";
ram(2641) <= "0000000000000000";
ram(2642) <= "0000000000000000";
ram(2643) <= "0000000000000000";
ram(2644) <= "0000000000000000";
ram(2645) <= "0000000000000000";
ram(2646) <= "0000000000000000";
ram(2647) <= "0000000000000000";
ram(2648) <= "0000000000000000";
ram(2649) <= "0000000000000000";
ram(2650) <= "0000000000000000";
ram(2651) <= "0000000000000000";
ram(2652) <= "0000000000000000";
ram(2653) <= "0000000000000000";
ram(2654) <= "0000000000000000";
ram(2655) <= "0000000000000000";
ram(2656) <= "0000000000000000";
ram(2657) <= "0000000000000000";
ram(2658) <= "0000000000000000";
ram(2659) <= "0000000000000000";
ram(2660) <= "0000000000000000";
ram(2661) <= "0000000000000000";
ram(2662) <= "0000000000000000";
ram(2663) <= "0000000000000000";
ram(2664) <= "0000000000000000";
ram(2665) <= "0000000000000000";
ram(2666) <= "0000000000000000";
ram(2667) <= "0000000000000000";
ram(2668) <= "0000000000000000";
ram(2669) <= "0000000000000000";
ram(2670) <= "0000000000000000";
ram(2671) <= "0000000000000000";
ram(2672) <= "0000000000000000";
ram(2673) <= "0000000000000000";
ram(2674) <= "0000000000000000";
ram(2675) <= "0000000000000000";
ram(2676) <= "0000000000000000";
ram(2677) <= "0000000000000000";
ram(2678) <= "0000000000000000";
ram(2679) <= "0000000000000000";
ram(2680) <= "0000000000000000";
ram(2681) <= "0000000000000000";
ram(2682) <= "0000000000000000";
ram(2683) <= "0000000000000000";
ram(2684) <= "0000000000000000";
ram(2685) <= "0000000000000000";
ram(2686) <= "0000000000000000";
ram(2687) <= "0000000000000000";
ram(2688) <= "0000000000000000";
ram(2689) <= "0000000000000000";
ram(2690) <= "0000000000000000";
ram(2691) <= "0000000000000000";
ram(2692) <= "0000000000000000";
ram(2693) <= "0000000000000000";
ram(2694) <= "0000000000000000";
ram(2695) <= "0000000000000000";
ram(2696) <= "0000000000000000";
ram(2697) <= "0000000000000000";
ram(2698) <= "0000000000000000";
ram(2699) <= "0000000000000000";
ram(2700) <= "0000000000000000";
ram(2701) <= "0000000000000000";
ram(2702) <= "0000000000000000";
ram(2703) <= "0000000000000000";
ram(2704) <= "0000000000000000";
ram(2705) <= "0000000000000000";
ram(2706) <= "0000000000000000";
ram(2707) <= "0000000000000000";
ram(2708) <= "0000000000000000";
ram(2709) <= "0000000000000000";
ram(2710) <= "0000000000000000";
ram(2711) <= "0000000000000000";
ram(2712) <= "0000000000000000";
ram(2713) <= "0000000000000000";
ram(2714) <= "0000000000000000";
ram(2715) <= "0000000000000000";
ram(2716) <= "0000000000000000";
ram(2717) <= "0000000000000000";
ram(2718) <= "0000000000000000";
ram(2719) <= "0000000000000000";
ram(2720) <= "0000000000000000";
ram(2721) <= "0000000000000000";
ram(2722) <= "0000000000000000";
ram(2723) <= "0000000000000000";
ram(2724) <= "0000000000000000";
ram(2725) <= "0000000000000000";
ram(2726) <= "0000000000000000";
ram(2727) <= "0000000000000000";
ram(2728) <= "0000000000000000";
ram(2729) <= "0000000000000000";
ram(2730) <= "0000000000000000";
ram(2731) <= "0000000000000000";
ram(2732) <= "0000000000000000";
ram(2733) <= "0000000000000000";
ram(2734) <= "0000000000000000";
ram(2735) <= "0000000000000000";
ram(2736) <= "0000000000000000";
ram(2737) <= "0000000000000000";
ram(2738) <= "0000000000000000";
ram(2739) <= "0000000000000000";
ram(2740) <= "0000000000000000";
ram(2741) <= "0000000000000000";
ram(2742) <= "0000000000000000";
ram(2743) <= "0000000000000000";
ram(2744) <= "0000000000000000";
ram(2745) <= "0000000000000000";
ram(2746) <= "0000000000000000";
ram(2747) <= "0000000000000000";
ram(2748) <= "0000000000000000";
ram(2749) <= "0000000000000000";
ram(2750) <= "0000000000000000";
ram(2751) <= "0000000000000000";
ram(2752) <= "0000000000000000";
ram(2753) <= "0000000000000000";
ram(2754) <= "0000000000000000";
ram(2755) <= "0000000000000000";
ram(2756) <= "0000000000000000";
ram(2757) <= "0000000000000000";
ram(2758) <= "0000000000000000";
ram(2759) <= "0000000000000000";
ram(2760) <= "0000000000000000";
ram(2761) <= "0000000000000000";
ram(2762) <= "0000000000000000";
ram(2763) <= "0000000000000000";
ram(2764) <= "0000000000000000";
ram(2765) <= "0000000000000000";
ram(2766) <= "0000000000000000";
ram(2767) <= "0000000000000000";
ram(2768) <= "0000000000000000";
ram(2769) <= "0000000000000000";
ram(2770) <= "0000000000000000";
ram(2771) <= "0000000000000000";
ram(2772) <= "0000000000000000";
ram(2773) <= "0000000000000000";
ram(2774) <= "0000000000000000";
ram(2775) <= "0000000000000000";
ram(2776) <= "0000000000000000";
ram(2777) <= "0000000000000000";
ram(2778) <= "0000000000000000";
ram(2779) <= "0000000000000000";
ram(2780) <= "0000000000000000";
ram(2781) <= "0000000000000000";
ram(2782) <= "0000000000000000";
ram(2783) <= "0000000000000000";
ram(2784) <= "0000000000000000";
ram(2785) <= "0000000000000000";
ram(2786) <= "0000000000000000";
ram(2787) <= "0000000000000000";
ram(2788) <= "0000000000000000";
ram(2789) <= "0000000000000000";
ram(2790) <= "0000000000000000";
ram(2791) <= "0000000000000000";
ram(2792) <= "0000000000000000";
ram(2793) <= "0000000000000000";
ram(2794) <= "0000000000000000";
ram(2795) <= "0000000000000000";
ram(2796) <= "0000000000000000";
ram(2797) <= "0000000000000000";
ram(2798) <= "0000000000000000";
ram(2799) <= "0000000000000000";
ram(2800) <= "0000000000000000";
ram(2801) <= "0000000000000000";
ram(2802) <= "0000000000000000";
ram(2803) <= "0000000000000000";
ram(2804) <= "0000000000000000";
ram(2805) <= "0000000000000000";
ram(2806) <= "0000000000000000";
ram(2807) <= "0000000000000000";
ram(2808) <= "0000000000000000";
ram(2809) <= "0000000000000000";
ram(2810) <= "0000000000000000";
ram(2811) <= "0000000000000000";
ram(2812) <= "0000000000000000";
ram(2813) <= "0000000000000000";
ram(2814) <= "0000000000000000";
ram(2815) <= "0000000000000000";
ram(2816) <= "0000000000000000";
ram(2817) <= "0000000000000000";
ram(2818) <= "0000000000000000";
ram(2819) <= "0000000000000000";
ram(2820) <= "0000000000000000";
ram(2821) <= "0000000000000000";
ram(2822) <= "0000000000000000";
ram(2823) <= "0000000000000000";
ram(2824) <= "0000000000000000";
ram(2825) <= "0000000000000000";
ram(2826) <= "0000000000000000";
ram(2827) <= "0000000000000000";
ram(2828) <= "0000000000000000";
ram(2829) <= "0000000000000000";
ram(2830) <= "0000000000000000";
ram(2831) <= "0000000000000000";
ram(2832) <= "0000000000000000";
ram(2833) <= "0000000000000000";
ram(2834) <= "0000000000000000";
ram(2835) <= "0000000000000000";
ram(2836) <= "0000000000000000";
ram(2837) <= "0000000000000000";
ram(2838) <= "0000000000000000";
ram(2839) <= "0000000000000000";
ram(2840) <= "0000000000000000";
ram(2841) <= "0000000000000000";
ram(2842) <= "0000000000000000";
ram(2843) <= "0000000000000000";
ram(2844) <= "0000000000000000";
ram(2845) <= "0000000000000000";
ram(2846) <= "0000000000000000";
ram(2847) <= "0000000000000000";
ram(2848) <= "0000000000000000";
ram(2849) <= "0000000000000000";
ram(2850) <= "0000000000000000";
ram(2851) <= "0000000000000000";
ram(2852) <= "0000000000000000";
ram(2853) <= "0000000000000000";
ram(2854) <= "0000000000000000";
ram(2855) <= "0000000000000000";
ram(2856) <= "0000000000000000";
ram(2857) <= "0000000000000000";
ram(2858) <= "0000000000000000";
ram(2859) <= "0000000000000000";
ram(2860) <= "0000000000000000";
ram(2861) <= "0000000000000000";
ram(2862) <= "0000000000000000";
ram(2863) <= "0000000000000000";
ram(2864) <= "0000000000000000";
ram(2865) <= "0000000000000000";
ram(2866) <= "0000000000000000";
ram(2867) <= "0000000000000000";
ram(2868) <= "0000000000000000";
ram(2869) <= "0000000000000000";
ram(2870) <= "0000000000000000";
ram(2871) <= "0000000000000000";
ram(2872) <= "0000000000000000";
ram(2873) <= "0000000000000000";
ram(2874) <= "0000000000000000";
ram(2875) <= "0000000000000000";
ram(2876) <= "0000000000000000";
ram(2877) <= "0000000000000000";
ram(2878) <= "0000000000000000";
ram(2879) <= "0000000000000000";
ram(2880) <= "0000000000000000";
ram(2881) <= "0000000000000000";
ram(2882) <= "0000000000000000";
ram(2883) <= "0000000000000000";
ram(2884) <= "0000000000000000";
ram(2885) <= "0000000000000000";
ram(2886) <= "0000000000000000";
ram(2887) <= "0000000000000000";
ram(2888) <= "0000000000000000";
ram(2889) <= "0000000000000000";
ram(2890) <= "0000000000000000";
ram(2891) <= "0000000000000000";
ram(2892) <= "0000000000000000";
ram(2893) <= "0000000000000000";
ram(2894) <= "0000000000000000";
ram(2895) <= "0000000000000000";
ram(2896) <= "0000000000000000";
ram(2897) <= "0000000000000000";
ram(2898) <= "0000000000000000";
ram(2899) <= "0000000000000000";
ram(2900) <= "0000000000000000";
ram(2901) <= "0000000000000000";
ram(2902) <= "0000000000000000";
ram(2903) <= "0000000000000000";
ram(2904) <= "0000000000000000";
ram(2905) <= "0000000000000000";
ram(2906) <= "0000000000000000";
ram(2907) <= "0000000000000000";
ram(2908) <= "0000000000000000";
ram(2909) <= "0000000000000000";
ram(2910) <= "0000000000000000";
ram(2911) <= "0000000000000000";
ram(2912) <= "0000000000000000";
ram(2913) <= "0000000000000000";
ram(2914) <= "0000000000000000";
ram(2915) <= "0000000000000000";
ram(2916) <= "0000000000000000";
ram(2917) <= "0000000000000000";
ram(2918) <= "0000000000000000";
ram(2919) <= "0000000000000000";
ram(2920) <= "0000000000000000";
ram(2921) <= "0000000000000000";
ram(2922) <= "0000000000000000";
ram(2923) <= "0000000000000000";
ram(2924) <= "0000000000000000";
ram(2925) <= "0000000000000000";
ram(2926) <= "0000000000000000";
ram(2927) <= "0000000000000000";
ram(2928) <= "0000000000000000";
ram(2929) <= "0000000000000000";
ram(2930) <= "0000000000000000";
ram(2931) <= "0000000000000000";
ram(2932) <= "0000000000000000";
ram(2933) <= "0000000000000000";
ram(2934) <= "0000000000000000";
ram(2935) <= "0000000000000000";
ram(2936) <= "0000000000000000";
ram(2937) <= "0000000000000000";
ram(2938) <= "0000000000000000";
ram(2939) <= "0000000000000000";
ram(2940) <= "0000000000000000";
ram(2941) <= "0000000000000000";
ram(2942) <= "0000000000000000";
ram(2943) <= "0000000000000000";
ram(2944) <= "0000000000000000";
ram(2945) <= "0000000000000000";
ram(2946) <= "0000000000000000";
ram(2947) <= "0000000000000000";
ram(2948) <= "0000000000000000";
ram(2949) <= "0000000000000000";
ram(2950) <= "0000000000000000";
ram(2951) <= "0000000000000000";
ram(2952) <= "0000000000000000";
ram(2953) <= "0000000000000000";
ram(2954) <= "0000000000000000";
ram(2955) <= "0000000000000000";
ram(2956) <= "0000000000000000";
ram(2957) <= "0000000000000000";
ram(2958) <= "0000000000000000";
ram(2959) <= "0000000000000000";
ram(2960) <= "0000000000000000";
ram(2961) <= "0000000000000000";
ram(2962) <= "0000000000000000";
ram(2963) <= "0000000000000000";
ram(2964) <= "0000000000000000";
ram(2965) <= "0000000000000000";
ram(2966) <= "0000000000000000";
ram(2967) <= "0000000000000000";
ram(2968) <= "0000000000000000";
ram(2969) <= "0000000000000000";
ram(2970) <= "0000000000000000";
ram(2971) <= "0000000000000000";
ram(2972) <= "0000000000000000";
ram(2973) <= "0000000000000000";
ram(2974) <= "0000000000000000";
ram(2975) <= "0000000000000000";
ram(2976) <= "0000000000000000";
ram(2977) <= "0000000000000000";
ram(2978) <= "0000000000000000";
ram(2979) <= "0000000000000000";
ram(2980) <= "0000000000000000";
ram(2981) <= "0000000000000000";
ram(2982) <= "0000000000000000";
ram(2983) <= "0000000000000000";
ram(2984) <= "0000000000000000";
ram(2985) <= "0000000000000000";
ram(2986) <= "0000000000000000";
ram(2987) <= "0000000000000000";
ram(2988) <= "0000000000000000";
ram(2989) <= "0000000000000000";
ram(2990) <= "0000000000000000";
ram(2991) <= "0000000000000000";
ram(2992) <= "0000000000000000";
ram(2993) <= "0000000000000000";
ram(2994) <= "0000000000000000";
ram(2995) <= "0000000000000000";
ram(2996) <= "0000000000000000";
ram(2997) <= "0000000000000000";
ram(2998) <= "0000000000000000";
ram(2999) <= "0000000000000000";
ram(3000) <= "0000000000000000";
ram(3001) <= "0000000000000000";
ram(3002) <= "0000000000000000";
ram(3003) <= "0000000000000000";
ram(3004) <= "0000000000000000";
ram(3005) <= "0000000000000000";
ram(3006) <= "0000000000000000";
ram(3007) <= "0000000000000000";
ram(3008) <= "0000000000000000";
ram(3009) <= "0000000000000000";
ram(3010) <= "0000000000000000";
ram(3011) <= "0000000000000000";
ram(3012) <= "0000000000000000";
ram(3013) <= "0000000000000000";
ram(3014) <= "0000000000000000";
ram(3015) <= "0000000000000000";
ram(3016) <= "0000000000000000";
ram(3017) <= "0000000000000000";
ram(3018) <= "0000000000000000";
ram(3019) <= "0000000000000000";
ram(3020) <= "0000000000000000";
ram(3021) <= "0000000000000000";
ram(3022) <= "0000000000000000";
ram(3023) <= "0000000000000000";
ram(3024) <= "0000000000000000";
ram(3025) <= "0000000000000000";
ram(3026) <= "0000000000000000";
ram(3027) <= "0000000000000000";
ram(3028) <= "0000000000000000";
ram(3029) <= "0000000000000000";
ram(3030) <= "0000000000000000";
ram(3031) <= "0000000000000000";
ram(3032) <= "0000000000000000";
ram(3033) <= "0000000000000000";
ram(3034) <= "0000000000000000";
ram(3035) <= "0000000000000000";
ram(3036) <= "0000000000000000";
ram(3037) <= "0000000000000000";
ram(3038) <= "0000000000000000";
ram(3039) <= "0000000000000000";
ram(3040) <= "0000000000000000";
ram(3041) <= "0000000000000000";
ram(3042) <= "0000000000000000";
ram(3043) <= "0000000000000000";
ram(3044) <= "0000000000000000";
ram(3045) <= "0000000000000000";
ram(3046) <= "0000000000000000";
ram(3047) <= "0000000000000000";
ram(3048) <= "0000000000000000";
ram(3049) <= "0000000000000000";
ram(3050) <= "0000000000000000";
ram(3051) <= "0000000000000000";
ram(3052) <= "0000000000000000";
ram(3053) <= "0000000000000000";
ram(3054) <= "0000000000000000";
ram(3055) <= "0000000000000000";
ram(3056) <= "0000000000000000";
ram(3057) <= "0000000000000000";
ram(3058) <= "0000000000000000";
ram(3059) <= "0000000000000000";
ram(3060) <= "0000000000000000";
ram(3061) <= "0000000000000000";
ram(3062) <= "0000000000000000";
ram(3063) <= "0000000000000000";
ram(3064) <= "0000000000000000";
ram(3065) <= "0000000000000000";
ram(3066) <= "0000000000000000";
ram(3067) <= "0000000000000000";
ram(3068) <= "0000000000000000";
ram(3069) <= "0000000000000000";
ram(3070) <= "0000000000000000";
ram(3071) <= "0000000000000000";
ram(3072) <= "0000000000000000";
ram(3073) <= "0000000000000000";
ram(3074) <= "0000000000000000";
ram(3075) <= "0000000000000000";
ram(3076) <= "0000000000000000";
ram(3077) <= "0000000000000000";
ram(3078) <= "0000000000000000";
ram(3079) <= "0000000000000000";
ram(3080) <= "0000000000000000";
ram(3081) <= "0000000000000000";
ram(3082) <= "0000000000000000";
ram(3083) <= "0000000000000000";
ram(3084) <= "0000000000000000";
ram(3085) <= "0000000000000000";
ram(3086) <= "0000000000000000";
ram(3087) <= "0000000000000000";
ram(3088) <= "0000000000000000";
ram(3089) <= "0000000000000000";
ram(3090) <= "0000000000000000";
ram(3091) <= "0000000000000000";
ram(3092) <= "0000000000000000";
ram(3093) <= "0000000000000000";
ram(3094) <= "0000000000000000";
ram(3095) <= "0000000000000000";
ram(3096) <= "0000000000000000";
ram(3097) <= "0000000000000000";
ram(3098) <= "0000000000000000";
ram(3099) <= "0000000000000000";
ram(3100) <= "0000000000000000";
ram(3101) <= "0000000000000000";
ram(3102) <= "0000000000000000";
ram(3103) <= "0000000000000000";
ram(3104) <= "0000000000000000";
ram(3105) <= "0000000000000000";
ram(3106) <= "0000000000000000";
ram(3107) <= "0000000000000000";
ram(3108) <= "0000000000000000";
ram(3109) <= "0000000000000000";
ram(3110) <= "0000000000000000";
ram(3111) <= "0000000000000000";
ram(3112) <= "0000000000000000";
ram(3113) <= "0000000000000000";
ram(3114) <= "0000000000000000";
ram(3115) <= "0000000000000000";
ram(3116) <= "0000000000000000";
ram(3117) <= "0000000000000000";
ram(3118) <= "0000000000000000";
ram(3119) <= "0000000000000000";
ram(3120) <= "0000000000000000";
ram(3121) <= "0000000000000000";
ram(3122) <= "0000000000000000";
ram(3123) <= "0000000000000000";
ram(3124) <= "0000000000000000";
ram(3125) <= "0000000000000000";
ram(3126) <= "0000000000000000";
ram(3127) <= "0000000000000000";
ram(3128) <= "0000000000000000";
ram(3129) <= "0000000000000000";
ram(3130) <= "0000000000000000";
ram(3131) <= "0000000000000000";
ram(3132) <= "0000000000000000";
ram(3133) <= "0000000000000000";
ram(3134) <= "0000000000000000";
ram(3135) <= "0000000000000000";
ram(3136) <= "0000000000000000";
ram(3137) <= "0000000000000000";
ram(3138) <= "0000000000000000";
ram(3139) <= "0000000000000000";
ram(3140) <= "0000000000000000";
ram(3141) <= "0000000000000000";
ram(3142) <= "0000000000000000";
ram(3143) <= "0000000000000000";
ram(3144) <= "0000000000000000";
ram(3145) <= "0000000000000000";
ram(3146) <= "0000000000000000";
ram(3147) <= "0000000000000000";
ram(3148) <= "0000000000000000";
ram(3149) <= "0000000000000000";
ram(3150) <= "0000000000000000";
ram(3151) <= "0000000000000000";
ram(3152) <= "0000000000000000";
ram(3153) <= "0000000000000000";
ram(3154) <= "0000000000000000";
ram(3155) <= "0000000000000000";
ram(3156) <= "0000000000000000";
ram(3157) <= "0000000000000000";
ram(3158) <= "0000000000000000";
ram(3159) <= "0000000000000000";
ram(3160) <= "0000000000000000";
ram(3161) <= "0000000000000000";
ram(3162) <= "0000000000000000";
ram(3163) <= "0000000000000000";
ram(3164) <= "0000000000000000";
ram(3165) <= "0000000000000000";
ram(3166) <= "0000000000000000";
ram(3167) <= "0000000000000000";
ram(3168) <= "0000000000000000";
ram(3169) <= "0000000000000000";
ram(3170) <= "0000000000000000";
ram(3171) <= "0000000000000000";
ram(3172) <= "0000000000000000";
ram(3173) <= "0000000000000000";
ram(3174) <= "0000000000000000";
ram(3175) <= "0000000000000000";
ram(3176) <= "0000000000000000";
ram(3177) <= "0000000000000000";
ram(3178) <= "0000000000000000";
ram(3179) <= "0000000000000000";
ram(3180) <= "0000000000000000";
ram(3181) <= "0000000000000000";
ram(3182) <= "0000000000000000";
ram(3183) <= "0000000000000000";
ram(3184) <= "0000000000000000";
ram(3185) <= "0000000000000000";
ram(3186) <= "0000000000000000";
ram(3187) <= "0000000000000000";
ram(3188) <= "0000000000000000";
ram(3189) <= "0000000000000000";
ram(3190) <= "0000000000000000";
ram(3191) <= "0000000000000000";
ram(3192) <= "0000000000000000";
ram(3193) <= "0000000000000000";
ram(3194) <= "0000000000000000";
ram(3195) <= "0000000000000000";
ram(3196) <= "0000000000000000";
ram(3197) <= "0000000000000000";
ram(3198) <= "0000000000000000";
ram(3199) <= "0000000000000000";
ram(3200) <= "0000000000000000";
ram(3201) <= "0000000000000000";
ram(3202) <= "0000000000000000";
ram(3203) <= "0000000000000000";
ram(3204) <= "0000000000000000";
ram(3205) <= "0000000000000000";
ram(3206) <= "0000000000000000";
ram(3207) <= "0000000000000000";
ram(3208) <= "0000000000000000";
ram(3209) <= "0000000000000000";
ram(3210) <= "0000000000000000";
ram(3211) <= "0000000000000000";
ram(3212) <= "0000000000000000";
ram(3213) <= "0000000000000000";
ram(3214) <= "0000000000000000";
ram(3215) <= "0000000000000000";
ram(3216) <= "0000000000000000";
ram(3217) <= "0000000000000000";
ram(3218) <= "0000000000000000";
ram(3219) <= "0000000000000000";
ram(3220) <= "0000000000000000";
ram(3221) <= "0000000000000000";
ram(3222) <= "0000000000000000";
ram(3223) <= "0000000000000000";
ram(3224) <= "0000000000000000";
ram(3225) <= "0000000000000000";
ram(3226) <= "0000000000000000";
ram(3227) <= "0000000000000000";
ram(3228) <= "0000000000000000";
ram(3229) <= "0000000000000000";
ram(3230) <= "0000000000000000";
ram(3231) <= "0000000000000000";
ram(3232) <= "0000000000000000";
ram(3233) <= "0000000000000000";
ram(3234) <= "0000000000000000";
ram(3235) <= "0000000000000000";
ram(3236) <= "0000000000000000";
ram(3237) <= "0000000000000000";
ram(3238) <= "0000000000000000";
ram(3239) <= "0000000000000000";
ram(3240) <= "0000000000000000";
ram(3241) <= "0000000000000000";
ram(3242) <= "0000000000000000";
ram(3243) <= "0000000000000000";
ram(3244) <= "0000000000000000";
ram(3245) <= "0000000000000000";
ram(3246) <= "0000000000000000";
ram(3247) <= "0000000000000000";
ram(3248) <= "0000000000000000";
ram(3249) <= "0000000000000000";
ram(3250) <= "0000000000000000";
ram(3251) <= "0000000000000000";
ram(3252) <= "0000000000000000";
ram(3253) <= "0000000000000000";
ram(3254) <= "0000000000000000";
ram(3255) <= "0000000000000000";
ram(3256) <= "0000000000000000";
ram(3257) <= "0000000000000000";
ram(3258) <= "0000000000000000";
ram(3259) <= "0000000000000000";
ram(3260) <= "0000000000000000";
ram(3261) <= "0000000000000000";
ram(3262) <= "0000000000000000";
ram(3263) <= "0000000000000000";
ram(3264) <= "0000000000000000";
ram(3265) <= "0000000000000000";
ram(3266) <= "0000000000000000";
ram(3267) <= "0000000000000000";
ram(3268) <= "0000000000000000";
ram(3269) <= "0000000000000000";
ram(3270) <= "0000000000000000";
ram(3271) <= "0000000000000000";
ram(3272) <= "0000000000000000";
ram(3273) <= "0000000000000000";
ram(3274) <= "0000000000000000";
ram(3275) <= "0000000000000000";
ram(3276) <= "0000000000000000";
ram(3277) <= "0000000000000000";
ram(3278) <= "0000000000000000";
ram(3279) <= "0000000000000000";
ram(3280) <= "0000000000000000";
ram(3281) <= "0000000000000000";
ram(3282) <= "0000000000000000";
ram(3283) <= "0000000000000000";
ram(3284) <= "0000000000000000";
ram(3285) <= "0000000000000000";
ram(3286) <= "0000000000000000";
ram(3287) <= "0000000000000000";
ram(3288) <= "0000000000000000";
ram(3289) <= "0000000000000000";
ram(3290) <= "0000000000000000";
ram(3291) <= "0000000000000000";
ram(3292) <= "0000000000000000";
ram(3293) <= "0000000000000000";
ram(3294) <= "0000000000000000";
ram(3295) <= "0000000000000000";
ram(3296) <= "0000000000000000";
ram(3297) <= "0000000000000000";
ram(3298) <= "0000000000000000";
ram(3299) <= "0000000000000000";
ram(3300) <= "0000000000000000";
ram(3301) <= "0000000000000000";
ram(3302) <= "0000000000000000";
ram(3303) <= "0000000000000000";
ram(3304) <= "0000000000000000";
ram(3305) <= "0000000000000000";
ram(3306) <= "0000000000000000";
ram(3307) <= "0000000000000000";
ram(3308) <= "0000000000000000";
ram(3309) <= "0000000000000000";
ram(3310) <= "0000000000000000";
ram(3311) <= "0000000000000000";
ram(3312) <= "0000000000000000";
ram(3313) <= "0000000000000000";
ram(3314) <= "0000000000000000";
ram(3315) <= "0000000000000000";
ram(3316) <= "0000000000000000";
ram(3317) <= "0000000000000000";
ram(3318) <= "0000000000000000";
ram(3319) <= "0000000000000000";
ram(3320) <= "0000000000000000";
ram(3321) <= "0000000000000000";
ram(3322) <= "0000000000000000";
ram(3323) <= "0000000000000000";
ram(3324) <= "0000000000000000";
ram(3325) <= "0000000000000000";
ram(3326) <= "0000000000000000";
ram(3327) <= "0000000000000000";
ram(3328) <= "0000000000000000";
ram(3329) <= "0000000000000000";
ram(3330) <= "0000000000000000";
ram(3331) <= "0000000000000000";
ram(3332) <= "0000000000000000";
ram(3333) <= "0000000000000000";
ram(3334) <= "0000000000000000";
ram(3335) <= "0000000000000000";
ram(3336) <= "0000000000000000";
ram(3337) <= "0000000000000000";
ram(3338) <= "0000000000000000";
ram(3339) <= "0000000000000000";
ram(3340) <= "0000000000000000";
ram(3341) <= "0000000000000000";
ram(3342) <= "0000000000000000";
ram(3343) <= "0000000000000000";
ram(3344) <= "0000000000000000";
ram(3345) <= "0000000000000000";
ram(3346) <= "0000000000000000";
ram(3347) <= "0000000000000000";
ram(3348) <= "0000000000000000";
ram(3349) <= "0000000000000000";
ram(3350) <= "0000000000000000";
ram(3351) <= "0000000000000000";
ram(3352) <= "0000000000000000";
ram(3353) <= "0000000000000000";
ram(3354) <= "0000000000000000";
ram(3355) <= "0000000000000000";
ram(3356) <= "0000000000000000";
ram(3357) <= "0000000000000000";
ram(3358) <= "0000000000000000";
ram(3359) <= "0000000000000000";
ram(3360) <= "0000000000000000";
ram(3361) <= "0000000000000000";
ram(3362) <= "0000000000000000";
ram(3363) <= "0000000000000000";
ram(3364) <= "0000000000000000";
ram(3365) <= "0000000000000000";
ram(3366) <= "0000000000000000";
ram(3367) <= "0000000000000000";
ram(3368) <= "0000000000000000";
ram(3369) <= "0000000000000000";
ram(3370) <= "0000000000000000";
ram(3371) <= "0000000000000000";
ram(3372) <= "0000000000000000";
ram(3373) <= "0000000000000000";
ram(3374) <= "0000000000000000";
ram(3375) <= "0000000000000000";
ram(3376) <= "0000000000000000";
ram(3377) <= "0000000000000000";
ram(3378) <= "0000000000000000";
ram(3379) <= "0000000000000000";
ram(3380) <= "0000000000000000";
ram(3381) <= "0000000000000000";
ram(3382) <= "0000000000000000";
ram(3383) <= "0000000000000000";
ram(3384) <= "0000000000000000";
ram(3385) <= "0000000000000000";
ram(3386) <= "0000000000000000";
ram(3387) <= "0000000000000000";
ram(3388) <= "0000000000000000";
ram(3389) <= "0000000000000000";
ram(3390) <= "0000000000000000";
ram(3391) <= "0000000000000000";
ram(3392) <= "0000000000000000";
ram(3393) <= "0000000000000000";
ram(3394) <= "0000000000000000";
ram(3395) <= "0000000000000000";
ram(3396) <= "0000000000000000";
ram(3397) <= "0000000000000000";
ram(3398) <= "0000000000000000";
ram(3399) <= "0000000000000000";
ram(3400) <= "0000000000000000";
ram(3401) <= "0000000000000000";
ram(3402) <= "0000000000000000";
ram(3403) <= "0000000000000000";
ram(3404) <= "0000000000000000";
ram(3405) <= "0000000000000000";
ram(3406) <= "0000000000000000";
ram(3407) <= "0000000000000000";
ram(3408) <= "0000000000000000";
ram(3409) <= "0000000000000000";
ram(3410) <= "0000000000000000";
ram(3411) <= "0000000000000000";
ram(3412) <= "0000000000000000";
ram(3413) <= "0000000000000000";
ram(3414) <= "0000000000000000";
ram(3415) <= "0000000000000000";
ram(3416) <= "0000000000000000";
ram(3417) <= "0000000000000000";
ram(3418) <= "0000000000000000";
ram(3419) <= "0000000000000000";
ram(3420) <= "0000000000000000";
ram(3421) <= "0000000000000000";
ram(3422) <= "0000000000000000";
ram(3423) <= "0000000000000000";
ram(3424) <= "0000000000000000";
ram(3425) <= "0000000000000000";
ram(3426) <= "0000000000000000";
ram(3427) <= "0000000000000000";
ram(3428) <= "0000000000000000";
ram(3429) <= "0000000000000000";
ram(3430) <= "0000000000000000";
ram(3431) <= "0000000000000000";
ram(3432) <= "0000000000000000";
ram(3433) <= "0000000000000000";
ram(3434) <= "0000000000000000";
ram(3435) <= "0000000000000000";
ram(3436) <= "0000000000000000";
ram(3437) <= "0000000000000000";
ram(3438) <= "0000000000000000";
ram(3439) <= "0000000000000000";
ram(3440) <= "0000000000000000";
ram(3441) <= "0000000000000000";
ram(3442) <= "0000000000000000";
ram(3443) <= "0000000000000000";
ram(3444) <= "0000000000000000";
ram(3445) <= "0000000000000000";
ram(3446) <= "0000000000000000";
ram(3447) <= "0000000000000000";
ram(3448) <= "0000000000000000";
ram(3449) <= "0000000000000000";
ram(3450) <= "0000000000000000";
ram(3451) <= "0000000000000000";
ram(3452) <= "0000000000000000";
ram(3453) <= "0000000000000000";
ram(3454) <= "0000000000000000";
ram(3455) <= "0000000000000000";
ram(3456) <= "0000000000000000";
ram(3457) <= "0000000000000000";
ram(3458) <= "0000000000000000";
ram(3459) <= "0000000000000000";
ram(3460) <= "0000000000000000";
ram(3461) <= "0000000000000000";
ram(3462) <= "0000000000000000";
ram(3463) <= "0000000000000000";
ram(3464) <= "0000000000000000";
ram(3465) <= "0000000000000000";
ram(3466) <= "0000000000000000";
ram(3467) <= "0000000000000000";
ram(3468) <= "0000000000000000";
ram(3469) <= "0000000000000000";
ram(3470) <= "0000000000000000";
ram(3471) <= "0000000000000000";
ram(3472) <= "0000000000000000";
ram(3473) <= "0000000000000000";
ram(3474) <= "0000000000000000";
ram(3475) <= "0000000000000000";
ram(3476) <= "0000000000000000";
ram(3477) <= "0000000000000000";
ram(3478) <= "0000000000000000";
ram(3479) <= "0000000000000000";
ram(3480) <= "0000000000000000";
ram(3481) <= "0000000000000000";
ram(3482) <= "0000000000000000";
ram(3483) <= "0000000000000000";
ram(3484) <= "0000000000000000";
ram(3485) <= "0000000000000000";
ram(3486) <= "0000000000000000";
ram(3487) <= "0000000000000000";
ram(3488) <= "0000000000000000";
ram(3489) <= "0000000000000000";
ram(3490) <= "0000000000000000";
ram(3491) <= "0000000000000000";
ram(3492) <= "0000000000000000";
ram(3493) <= "0000000000000000";
ram(3494) <= "0000000000000000";
ram(3495) <= "0000000000000000";
ram(3496) <= "0000000000000000";
ram(3497) <= "0000000000000000";
ram(3498) <= "0000000000000000";
ram(3499) <= "0000000000000000";
ram(3500) <= "0000000000000000";
ram(3501) <= "0000000000000000";
ram(3502) <= "0000000000000000";
ram(3503) <= "0000000000000000";
ram(3504) <= "0000000000000000";
ram(3505) <= "0000000000000000";
ram(3506) <= "0000000000000000";
ram(3507) <= "0000000000000000";
ram(3508) <= "0000000000000000";
ram(3509) <= "0000000000000000";
ram(3510) <= "0000000000000000";
ram(3511) <= "0000000000000000";
ram(3512) <= "0000000000000000";
ram(3513) <= "0000000000000000";
ram(3514) <= "0000000000000000";
ram(3515) <= "0000000000000000";
ram(3516) <= "0000000000000000";
ram(3517) <= "0000000000000000";
ram(3518) <= "0000000000000000";
ram(3519) <= "0000000000000000";
ram(3520) <= "0000000000000000";
ram(3521) <= "0000000000000000";
ram(3522) <= "0000000000000000";
ram(3523) <= "0000000000000000";
ram(3524) <= "0000000000000000";
ram(3525) <= "0000000000000000";
ram(3526) <= "0000000000000000";
ram(3527) <= "0000000000000000";
ram(3528) <= "0000000000000000";
ram(3529) <= "0000000000000000";
ram(3530) <= "0000000000000000";
ram(3531) <= "0000000000000000";
ram(3532) <= "0000000000000000";
ram(3533) <= "0000000000000000";
ram(3534) <= "0000000000000000";
ram(3535) <= "0000000000000000";
ram(3536) <= "0000000000000000";
ram(3537) <= "0000000000000000";
ram(3538) <= "0000000000000000";
ram(3539) <= "0000000000000000";
ram(3540) <= "0000000000000000";
ram(3541) <= "0000000000000000";
ram(3542) <= "0000000000000000";
ram(3543) <= "0000000000000000";
ram(3544) <= "0000000000000000";
ram(3545) <= "0000000000000000";
ram(3546) <= "0000000000000000";
ram(3547) <= "0000000000000000";
ram(3548) <= "0000000000000000";
ram(3549) <= "0000000000000000";
ram(3550) <= "0000000000000000";
ram(3551) <= "0000000000000000";
ram(3552) <= "0000000000000000";
ram(3553) <= "0000000000000000";
ram(3554) <= "0000000000000000";
ram(3555) <= "0000000000000000";
ram(3556) <= "0000000000000000";
ram(3557) <= "0000000000000000";
ram(3558) <= "0000000000000000";
ram(3559) <= "0000000000000000";
ram(3560) <= "0000000000000000";
ram(3561) <= "0000000000000000";
ram(3562) <= "0000000000000000";
ram(3563) <= "0000000000000000";
ram(3564) <= "0000000000000000";
ram(3565) <= "0000000000000000";
ram(3566) <= "0000000000000000";
ram(3567) <= "0000000000000000";
ram(3568) <= "0000000000000000";
ram(3569) <= "0000000000000000";
ram(3570) <= "0000000000000000";
ram(3571) <= "0000000000000000";
ram(3572) <= "0000000000000000";
ram(3573) <= "0000000000000000";
ram(3574) <= "0000000000000000";
ram(3575) <= "0000000000000000";
ram(3576) <= "0000000000000000";
ram(3577) <= "0000000000000000";
ram(3578) <= "0000000000000000";
ram(3579) <= "0000000000000000";
ram(3580) <= "0000000000000000";
ram(3581) <= "0000000000000000";
ram(3582) <= "0000000000000000";
ram(3583) <= "0000000000000000";
ram(3584) <= "0000000000000000";
ram(3585) <= "0000000000000000";
ram(3586) <= "0000000000000000";
ram(3587) <= "0000000000000000";
ram(3588) <= "0000000000000000";
ram(3589) <= "0000000000000000";
ram(3590) <= "0000000000000000";
ram(3591) <= "0000000000000000";
ram(3592) <= "0000000000000000";
ram(3593) <= "0000000000000000";
ram(3594) <= "0000000000000000";
ram(3595) <= "0000000000000000";
ram(3596) <= "0000000000000000";
ram(3597) <= "0000000000000000";
ram(3598) <= "0000000000000000";
ram(3599) <= "0000000000000000";
ram(3600) <= "0000000000000000";
ram(3601) <= "0000000000000000";
ram(3602) <= "0000000000000000";
ram(3603) <= "0000000000000000";
ram(3604) <= "0000000000000000";
ram(3605) <= "0000000000000000";
ram(3606) <= "0000000000000000";
ram(3607) <= "0000000000000000";
ram(3608) <= "0000000000000000";
ram(3609) <= "0000000000000000";
ram(3610) <= "0000000000000000";
ram(3611) <= "0000000000000000";
ram(3612) <= "0000000000000000";
ram(3613) <= "0000000000000000";
ram(3614) <= "0000000000000000";
ram(3615) <= "0000000000000000";
ram(3616) <= "0000000000000000";
ram(3617) <= "0000000000000000";
ram(3618) <= "0000000000000000";
ram(3619) <= "0000000000000000";
ram(3620) <= "0000000000000000";
ram(3621) <= "0000000000000000";
ram(3622) <= "0000000000000000";
ram(3623) <= "0000000000000000";
ram(3624) <= "0000000000000000";
ram(3625) <= "0000000000000000";
ram(3626) <= "0000000000000000";
ram(3627) <= "0000000000000000";
ram(3628) <= "0000000000000000";
ram(3629) <= "0000000000000000";
ram(3630) <= "0000000000000000";
ram(3631) <= "0000000000000000";
ram(3632) <= "0000000000000000";
ram(3633) <= "0000000000000000";
ram(3634) <= "0000000000000000";
ram(3635) <= "0000000000000000";
ram(3636) <= "0000000000000000";
ram(3637) <= "0000000000000000";
ram(3638) <= "0000000000000000";
ram(3639) <= "0000000000000000";
ram(3640) <= "0000000000000000";
ram(3641) <= "0000000000000000";
ram(3642) <= "0000000000000000";
ram(3643) <= "0000000000000000";
ram(3644) <= "0000000000000000";
ram(3645) <= "0000000000000000";
ram(3646) <= "0000000000000000";
ram(3647) <= "0000000000000000";
ram(3648) <= "0000000000000000";
ram(3649) <= "0000000000000000";
ram(3650) <= "0000000000000000";
ram(3651) <= "0000000000000000";
ram(3652) <= "0000000000000000";
ram(3653) <= "0000000000000000";
ram(3654) <= "0000000000000000";
ram(3655) <= "0000000000000000";
ram(3656) <= "0000000000000000";
ram(3657) <= "0000000000000000";
ram(3658) <= "0000000000000000";
ram(3659) <= "0000000000000000";
ram(3660) <= "0000000000000000";
ram(3661) <= "0000000000000000";
ram(3662) <= "0000000000000000";
ram(3663) <= "0000000000000000";
ram(3664) <= "0000000000000000";
ram(3665) <= "0000000000000000";
ram(3666) <= "0000000000000000";
ram(3667) <= "0000000000000000";
ram(3668) <= "0000000000000000";
ram(3669) <= "0000000000000000";
ram(3670) <= "0000000000000000";
ram(3671) <= "0000000000000000";
ram(3672) <= "0000000000000000";
ram(3673) <= "0000000000000000";
ram(3674) <= "0000000000000000";
ram(3675) <= "0000000000000000";
ram(3676) <= "0000000000000000";
ram(3677) <= "0000000000000000";
ram(3678) <= "0000000000000000";
ram(3679) <= "0000000000000000";
ram(3680) <= "0000000000000000";
ram(3681) <= "0000000000000000";
ram(3682) <= "0000000000000000";
ram(3683) <= "0000000000000000";
ram(3684) <= "0000000000000000";
ram(3685) <= "0000000000000000";
ram(3686) <= "0000000000000000";
ram(3687) <= "0000000000000000";
ram(3688) <= "0000000000000000";
ram(3689) <= "0000000000000000";
ram(3690) <= "0000000000000000";
ram(3691) <= "0000000000000000";
ram(3692) <= "0000000000000000";
ram(3693) <= "0000000000000000";
ram(3694) <= "0000000000000000";
ram(3695) <= "0000000000000000";
ram(3696) <= "0000000000000000";
ram(3697) <= "0000000000000000";
ram(3698) <= "0000000000000000";
ram(3699) <= "0000000000000000";
ram(3700) <= "0000000000000000";
ram(3701) <= "0000000000000000";
ram(3702) <= "0000000000000000";
ram(3703) <= "0000000000000000";
ram(3704) <= "0000000000000000";
ram(3705) <= "0000000000000000";
ram(3706) <= "0000000000000000";
ram(3707) <= "0000000000000000";
ram(3708) <= "0000000000000000";
ram(3709) <= "0000000000000000";
ram(3710) <= "0000000000000000";
ram(3711) <= "0000000000000000";
ram(3712) <= "0000000000000000";
ram(3713) <= "0000000000000000";
ram(3714) <= "0000000000000000";
ram(3715) <= "0000000000000000";
ram(3716) <= "0000000000000000";
ram(3717) <= "0000000000000000";
ram(3718) <= "0000000000000000";
ram(3719) <= "0000000000000000";
ram(3720) <= "0000000000000000";
ram(3721) <= "0000000000000000";
ram(3722) <= "0000000000000000";
ram(3723) <= "0000000000000000";
ram(3724) <= "0000000000000000";
ram(3725) <= "0000000000000000";
ram(3726) <= "0000000000000000";
ram(3727) <= "0000000000000000";
ram(3728) <= "0000000000000000";
ram(3729) <= "0000000000000000";
ram(3730) <= "0000000000000000";
ram(3731) <= "0000000000000000";
ram(3732) <= "0000000000000000";
ram(3733) <= "0000000000000000";
ram(3734) <= "0000000000000000";
ram(3735) <= "0000000000000000";
ram(3736) <= "0000000000000000";
ram(3737) <= "0000000000000000";
ram(3738) <= "0000000000000000";
ram(3739) <= "0000000000000000";
ram(3740) <= "0000000000000000";
ram(3741) <= "0000000000000000";
ram(3742) <= "0000000000000000";
ram(3743) <= "0000000000000000";
ram(3744) <= "0000000000000000";
ram(3745) <= "0000000000000000";
ram(3746) <= "0000000000000000";
ram(3747) <= "0000000000000000";
ram(3748) <= "0000000000000000";
ram(3749) <= "0000000000000000";
ram(3750) <= "0000000000000000";
ram(3751) <= "0000000000000000";
ram(3752) <= "0000000000000000";
ram(3753) <= "0000000000000000";
ram(3754) <= "0000000000000000";
ram(3755) <= "0000000000000000";
ram(3756) <= "0000000000000000";
ram(3757) <= "0000000000000000";
ram(3758) <= "0000000000000000";
ram(3759) <= "0000000000000000";
ram(3760) <= "0000000000000000";
ram(3761) <= "0000000000000000";
ram(3762) <= "0000000000000000";
ram(3763) <= "0000000000000000";
ram(3764) <= "0000000000000000";
ram(3765) <= "0000000000000000";
ram(3766) <= "0000000000000000";
ram(3767) <= "0000000000000000";
ram(3768) <= "0000000000000000";
ram(3769) <= "0000000000000000";
ram(3770) <= "0000000000000000";
ram(3771) <= "0000000000000000";
ram(3772) <= "0000000000000000";
ram(3773) <= "0000000000000000";
ram(3774) <= "0000000000000000";
ram(3775) <= "0000000000000000";
ram(3776) <= "0000000000000000";
ram(3777) <= "0000000000000000";
ram(3778) <= "0000000000000000";
ram(3779) <= "0000000000000000";
ram(3780) <= "0000000000000000";
ram(3781) <= "0000000000000000";
ram(3782) <= "0000000000000000";
ram(3783) <= "0000000000000000";
ram(3784) <= "0000000000000000";
ram(3785) <= "0000000000000000";
ram(3786) <= "0000000000000000";
ram(3787) <= "0000000000000000";
ram(3788) <= "0000000000000000";
ram(3789) <= "0000000000000000";
ram(3790) <= "0000000000000000";
ram(3791) <= "0000000000000000";
ram(3792) <= "0000000000000000";
ram(3793) <= "0000000000000000";
ram(3794) <= "0000000000000000";
ram(3795) <= "0000000000000000";
ram(3796) <= "0000000000000000";
ram(3797) <= "0000000000000000";
ram(3798) <= "0000000000000000";
ram(3799) <= "0000000000000000";
ram(3800) <= "0000000000000000";
ram(3801) <= "0000000000000000";
ram(3802) <= "0000000000000000";
ram(3803) <= "0000000000000000";
ram(3804) <= "0000000000000000";
ram(3805) <= "0000000000000000";
ram(3806) <= "0000000000000000";
ram(3807) <= "0000000000000000";
ram(3808) <= "0000000000000000";
ram(3809) <= "0000000000000000";
ram(3810) <= "0000000000000000";
ram(3811) <= "0000000000000000";
ram(3812) <= "0000000000000000";
ram(3813) <= "0000000000000000";
ram(3814) <= "0000000000000000";
ram(3815) <= "0000000000000000";
ram(3816) <= "0000000000000000";
ram(3817) <= "0000000000000000";
ram(3818) <= "0000000000000000";
ram(3819) <= "0000000000000000";
ram(3820) <= "0000000000000000";
ram(3821) <= "0000000000000000";
ram(3822) <= "0000000000000000";
ram(3823) <= "0000000000000000";
ram(3824) <= "0000000000000000";
ram(3825) <= "0000000000000000";
ram(3826) <= "0000000000000000";
ram(3827) <= "0000000000000000";
ram(3828) <= "0000000000000000";
ram(3829) <= "0000000000000000";
ram(3830) <= "0000000000000000";
ram(3831) <= "0000000000000000";
ram(3832) <= "0000000000000000";
ram(3833) <= "0000000000000000";
ram(3834) <= "0000000000000000";
ram(3835) <= "0000000000000000";
ram(3836) <= "0000000000000000";
ram(3837) <= "0000000000000000";
ram(3838) <= "0000000000000000";
ram(3839) <= "0000000000000000";
ram(3840) <= "0000000000000000";
ram(3841) <= "0000000000000000";
ram(3842) <= "0000000000000000";
ram(3843) <= "0000000000000000";
ram(3844) <= "0000000000000000";
ram(3845) <= "0000000000000000";
ram(3846) <= "0000000000000000";
ram(3847) <= "0000000000000000";
ram(3848) <= "0000000000000000";
ram(3849) <= "0000000000000000";
ram(3850) <= "0000000000000000";
ram(3851) <= "0000000000000000";
ram(3852) <= "0000000000000000";
ram(3853) <= "0000000000000000";
ram(3854) <= "0000000000000000";
ram(3855) <= "0000000000000000";
ram(3856) <= "0000000000000000";
ram(3857) <= "0000000000000000";
ram(3858) <= "0000000000000000";
ram(3859) <= "0000000000000000";
ram(3860) <= "0000000000000000";
ram(3861) <= "0000000000000000";
ram(3862) <= "0000000000000000";
ram(3863) <= "0000000000000000";
ram(3864) <= "0000000000000000";
ram(3865) <= "0000000000000000";
ram(3866) <= "0000000000000000";
ram(3867) <= "0000000000000000";
ram(3868) <= "0000000000000000";
ram(3869) <= "0000000000000000";
ram(3870) <= "0000000000000000";
ram(3871) <= "0000000000000000";
ram(3872) <= "0000000000000000";
ram(3873) <= "0000000000000000";
ram(3874) <= "0000000000000000";
ram(3875) <= "0000000000000000";
ram(3876) <= "0000000000000000";
ram(3877) <= "0000000000000000";
ram(3878) <= "0000000000000000";
ram(3879) <= "0000000000000000";
ram(3880) <= "0000000000000000";
ram(3881) <= "0000000000000000";
ram(3882) <= "0000000000000000";
ram(3883) <= "0000000000000000";
ram(3884) <= "0000000000000000";
ram(3885) <= "0000000000000000";
ram(3886) <= "0000000000000000";
ram(3887) <= "0000000000000000";
ram(3888) <= "0000000000000000";
ram(3889) <= "0000000000000000";
ram(3890) <= "0000000000000000";
ram(3891) <= "0000000000000000";
ram(3892) <= "0000000000000000";
ram(3893) <= "0000000000000000";
ram(3894) <= "0000000000000000";
ram(3895) <= "0000000000000000";
ram(3896) <= "0000000000000000";
ram(3897) <= "0000000000000000";
ram(3898) <= "0000000000000000";
ram(3899) <= "0000000000000000";
ram(3900) <= "0000000000000000";
ram(3901) <= "0000000000000000";
ram(3902) <= "0000000000000000";
ram(3903) <= "0000000000000000";
ram(3904) <= "0000000000000000";
ram(3905) <= "0000000000000000";
ram(3906) <= "0000000000000000";
ram(3907) <= "0000000000000000";
ram(3908) <= "0000000000000000";
ram(3909) <= "0000000000000000";
ram(3910) <= "0000000000000000";
ram(3911) <= "0000000000000000";
ram(3912) <= "0000000000000000";
ram(3913) <= "0000000000000000";
ram(3914) <= "0000000000000000";
ram(3915) <= "0000000000000000";
ram(3916) <= "0000000000000000";
ram(3917) <= "0000000000000000";
ram(3918) <= "0000000000000000";
ram(3919) <= "0000000000000000";
ram(3920) <= "0000000000000000";
ram(3921) <= "0000000000000000";
ram(3922) <= "0000000000000000";
ram(3923) <= "0000000000000000";
ram(3924) <= "0000000000000000";
ram(3925) <= "0000000000000000";
ram(3926) <= "0000000000000000";
ram(3927) <= "0000000000000000";
ram(3928) <= "0000000000000000";
ram(3929) <= "0000000000000000";
ram(3930) <= "0000000000000000";
ram(3931) <= "0000000000000000";
ram(3932) <= "0000000000000000";
ram(3933) <= "0000000000000000";
ram(3934) <= "0000000000000000";
ram(3935) <= "0000000000000000";
ram(3936) <= "0000000000000000";
ram(3937) <= "0000000000000000";
ram(3938) <= "0000000000000000";
ram(3939) <= "0000000000000000";
ram(3940) <= "0000000000000000";
ram(3941) <= "0000000000000000";
ram(3942) <= "0000000000000000";
ram(3943) <= "0000000000000000";
ram(3944) <= "0000000000000000";
ram(3945) <= "0000000000000000";
ram(3946) <= "0000000000000000";
ram(3947) <= "0000000000000000";
ram(3948) <= "0000000000000000";
ram(3949) <= "0000000000000000";
ram(3950) <= "0000000000000000";
ram(3951) <= "0000000000000000";
ram(3952) <= "0000000000000000";
ram(3953) <= "0000000000000000";
ram(3954) <= "0000000000000000";
ram(3955) <= "0000000000000000";
ram(3956) <= "0000000000000000";
ram(3957) <= "0000000000000000";
ram(3958) <= "0000000000000000";
ram(3959) <= "0000000000000000";
ram(3960) <= "0000000000000000";
ram(3961) <= "0000000000000000";
ram(3962) <= "0000000000000000";
ram(3963) <= "0000000000000000";
ram(3964) <= "0000000000000000";
ram(3965) <= "0000000000000000";
ram(3966) <= "0000000000000000";
ram(3967) <= "0000000000000000";
ram(3968) <= "0000000000000000";
ram(3969) <= "0000000000000000";
ram(3970) <= "0000000000000000";
ram(3971) <= "0000000000000000";
ram(3972) <= "0000000000000000";
ram(3973) <= "0000000000000000";
ram(3974) <= "0000000000000000";
ram(3975) <= "0000000000000000";
ram(3976) <= "0000000000000000";
ram(3977) <= "0000000000000000";
ram(3978) <= "0000000000000000";
ram(3979) <= "0000000000000000";
ram(3980) <= "0000000000000000";
ram(3981) <= "0000000000000000";
ram(3982) <= "0000000000000000";
ram(3983) <= "0000000000000000";
ram(3984) <= "0000000000000000";
ram(3985) <= "0000000000000000";
ram(3986) <= "0000000000000000";
ram(3987) <= "0000000000000000";
ram(3988) <= "0000000000000000";
ram(3989) <= "0000000000000000";
ram(3990) <= "0000000000000000";
ram(3991) <= "0000000000000000";
ram(3992) <= "0000000000000000";
ram(3993) <= "0000000000000000";
ram(3994) <= "0000000000000000";
ram(3995) <= "0000000000000000";
ram(3996) <= "0000000000000000";
ram(3997) <= "0000000000000000";
ram(3998) <= "0000000000000000";
ram(3999) <= "0000000000000000";
ram(4000) <= "0000000000000000";
ram(4001) <= "0000000000000000";
ram(4002) <= "0000000000000000";
ram(4003) <= "0000000000000000";
ram(4004) <= "0000000000000000";
ram(4005) <= "0000000000000000";
ram(4006) <= "0000000000000000";
ram(4007) <= "0000000000000000";
ram(4008) <= "0000000000000000";
ram(4009) <= "0000000000000000";
ram(4010) <= "0000000000000000";
ram(4011) <= "0000000000000000";
ram(4012) <= "0000000000000000";
ram(4013) <= "0000000000000000";
ram(4014) <= "0000000000000000";
ram(4015) <= "0000000000000000";
ram(4016) <= "0000000000000000";
ram(4017) <= "0000000000000000";
ram(4018) <= "0000000000000000";
ram(4019) <= "0000000000000000";
ram(4020) <= "0000000000000000";
ram(4021) <= "0000000000000000";
ram(4022) <= "0000000000000000";
ram(4023) <= "0000000000000000";
ram(4024) <= "0000000000000000";
ram(4025) <= "0000000000000000";
ram(4026) <= "0000000000000000";
ram(4027) <= "0000000000000000";
ram(4028) <= "0000000000000000";
ram(4029) <= "0000000000000000";
ram(4030) <= "0000000000000000";
ram(4031) <= "0000000000000000";
ram(4032) <= "0000000000000000";
ram(4033) <= "0000000000000000";
ram(4034) <= "0000000000000000";
ram(4035) <= "0000000000000000";
ram(4036) <= "0000000000000000";
ram(4037) <= "0000000000000000";
ram(4038) <= "0000000000000000";
ram(4039) <= "0000000000000000";
ram(4040) <= "0000000000000000";
ram(4041) <= "0000000000000000";
ram(4042) <= "0000000000000000";
ram(4043) <= "0000000000000000";
ram(4044) <= "0000000000000000";
ram(4045) <= "0000000000000000";
ram(4046) <= "0000000000000000";
ram(4047) <= "0000000000000000";
ram(4048) <= "0000000000000000";
ram(4049) <= "0000000000000000";
ram(4050) <= "0000000000000000";
ram(4051) <= "0000000000000000";
ram(4052) <= "0000000000000000";
ram(4053) <= "0000000000000000";
ram(4054) <= "0000000000000000";
ram(4055) <= "0000000000000000";
ram(4056) <= "0000000000000000";
ram(4057) <= "0000000000000000";
ram(4058) <= "0000000000000000";
ram(4059) <= "0000000000000000";
ram(4060) <= "0000000000000000";
ram(4061) <= "0000000000000000";
ram(4062) <= "0000000000000000";
ram(4063) <= "0000000000000000";
ram(4064) <= "0000000000000000";
ram(4065) <= "0000000000000000";
ram(4066) <= "0000000000000000";
ram(4067) <= "0000000000000000";
ram(4068) <= "0000000000000000";
ram(4069) <= "0000000000000000";
ram(4070) <= "0000000000000000";
ram(4071) <= "0000000000000000";
ram(4072) <= "0000000000000000";
ram(4073) <= "0000000000000000";
ram(4074) <= "0000000000000000";
ram(4075) <= "0000000000000000";
ram(4076) <= "0000000000000000";
ram(4077) <= "0000000000000000";
ram(4078) <= "0000000000000000";
ram(4079) <= "0000000000000000";
ram(4080) <= "0000000000000000";
ram(4081) <= "0000000000000000";
ram(4082) <= "0000000000000000";
ram(4083) <= "0000000000000000";
ram(4084) <= "0000000000000000";
ram(4085) <= "0000000000000000";
ram(4086) <= "0000000000000000";
ram(4087) <= "0000000000000000";
ram(4088) <= "0000000000000000";
ram(4089) <= "0000000000000000";
ram(4090) <= "0000000000000000";
ram(4091) <= "0000000000000000";
ram(4092) <= "0000000000000000";
ram(4093) <= "0000000000000000";
ram(4094) <= "0000000000000000";
ram(4095) <= "0000000000000000";
